module fetch_unit_DW01_add_0 (
	A, 
	B, 
	CI, 
	SUM, 
	CO);
   input [31:0] A;
   input [31:0] B;
   input CI;
   output [31:0] SUM;
   output CO;

   // Internal wires
   wire n30;
   wire n31;
   wire n32;
   wire n33;
   wire n34;
   wire n35;
   wire n36;
   wire n37;
   wire n38;
   wire n39;
   wire n40;
   wire n41;
   wire n42;
   wire n43;
   wire n44;
   wire n45;
   wire n46;
   wire n47;
   wire n48;
   wire n49;
   wire n50;
   wire n51;
   wire n52;
   wire n53;
   wire n54;
   wire n55;
   wire n56;
   wire n57;

   assign SUM[1] = A[1] ;
   assign SUM[0] = A[0] ;

   XOR2_X1 U1 (.A(A[20]),
	.B(n43),
	.Z(SUM[20]));
   XOR2_X1 U2 (.A(A[19]),
	.B(n44),
	.Z(SUM[19]));
   XOR2_X1 U3 (.A(A[18]),
	.B(n45),
	.Z(SUM[18]));
   XOR2_X1 U4 (.A(A[17]),
	.B(n46),
	.Z(SUM[17]));
   XNOR2_X1 U5 (.A(A[31]),
	.B(n57),
	.ZN(SUM[31]));
   XOR2_X1 U6 (.A(A[3]),
	.B(A[2]),
	.Z(SUM[3]));
   XOR2_X1 U7 (.A(A[16]),
	.B(n47),
	.Z(SUM[16]));
   XOR2_X1 U8 (.A(A[15]),
	.B(n48),
	.Z(SUM[15]));
   XOR2_X1 U9 (.A(A[14]),
	.B(n49),
	.Z(SUM[14]));
   XOR2_X1 U10 (.A(A[13]),
	.B(n50),
	.Z(SUM[13]));
   XOR2_X1 U11 (.A(A[12]),
	.B(n51),
	.Z(SUM[12]));
   XOR2_X1 U12 (.A(A[11]),
	.B(n52),
	.Z(SUM[11]));
   XOR2_X1 U13 (.A(A[10]),
	.B(n53),
	.Z(SUM[10]));
   XOR2_X1 U14 (.A(A[9]),
	.B(n54),
	.Z(SUM[9]));
   XOR2_X1 U15 (.A(A[8]),
	.B(n55),
	.Z(SUM[8]));
   XOR2_X1 U16 (.A(A[7]),
	.B(n30),
	.Z(SUM[7]));
   XOR2_X1 U17 (.A(A[6]),
	.B(n31),
	.Z(SUM[6]));
   XOR2_X1 U18 (.A(A[5]),
	.B(n32),
	.Z(SUM[5]));
   XOR2_X1 U19 (.A(A[4]),
	.B(n56),
	.Z(SUM[4]));
   XOR2_X1 U20 (.A(A[23]),
	.B(n40),
	.Z(SUM[23]));
   XOR2_X1 U21 (.A(A[22]),
	.B(n41),
	.Z(SUM[22]));
   XOR2_X1 U22 (.A(A[21]),
	.B(n42),
	.Z(SUM[21]));
   XOR2_X1 U23 (.A(A[30]),
	.B(n33),
	.Z(SUM[30]));
   XOR2_X1 U24 (.A(A[29]),
	.B(n34),
	.Z(SUM[29]));
   XOR2_X1 U25 (.A(A[28]),
	.B(n35),
	.Z(SUM[28]));
   XOR2_X1 U26 (.A(A[27]),
	.B(n36),
	.Z(SUM[27]));
   XOR2_X1 U27 (.A(A[26]),
	.B(n37),
	.Z(SUM[26]));
   XOR2_X1 U28 (.A(A[24]),
	.B(n39),
	.Z(SUM[24]));
   XOR2_X1 U29 (.A(A[25]),
	.B(n38),
	.Z(SUM[25]));
   NAND2_X1 U30 (.A1(A[30]),
	.A2(n33),
	.ZN(n57));
   AND2_X1 U31 (.A1(A[6]),
	.A2(n31),
	.ZN(n30));
   AND2_X1 U32 (.A1(A[5]),
	.A2(n32),
	.ZN(n31));
   AND2_X1 U33 (.A1(A[4]),
	.A2(n56),
	.ZN(n32));
   AND2_X1 U34 (.A1(A[29]),
	.A2(n34),
	.ZN(n33));
   AND2_X1 U35 (.A1(A[28]),
	.A2(n35),
	.ZN(n34));
   AND2_X1 U36 (.A1(A[27]),
	.A2(n36),
	.ZN(n35));
   AND2_X1 U37 (.A1(A[26]),
	.A2(n37),
	.ZN(n36));
   AND2_X1 U38 (.A1(A[25]),
	.A2(n38),
	.ZN(n37));
   AND2_X1 U39 (.A1(A[24]),
	.A2(n39),
	.ZN(n38));
   AND2_X1 U40 (.A1(A[23]),
	.A2(n40),
	.ZN(n39));
   AND2_X1 U41 (.A1(A[22]),
	.A2(n41),
	.ZN(n40));
   AND2_X1 U42 (.A1(A[21]),
	.A2(n42),
	.ZN(n41));
   AND2_X1 U43 (.A1(A[20]),
	.A2(n43),
	.ZN(n42));
   AND2_X1 U44 (.A1(A[19]),
	.A2(n44),
	.ZN(n43));
   AND2_X1 U45 (.A1(A[18]),
	.A2(n45),
	.ZN(n44));
   AND2_X1 U46 (.A1(A[17]),
	.A2(n46),
	.ZN(n45));
   AND2_X1 U47 (.A1(A[16]),
	.A2(n47),
	.ZN(n46));
   AND2_X1 U48 (.A1(A[15]),
	.A2(n48),
	.ZN(n47));
   AND2_X1 U49 (.A1(A[14]),
	.A2(n49),
	.ZN(n48));
   AND2_X1 U50 (.A1(A[13]),
	.A2(n50),
	.ZN(n49));
   AND2_X1 U51 (.A1(A[12]),
	.A2(n51),
	.ZN(n50));
   AND2_X1 U52 (.A1(A[11]),
	.A2(n52),
	.ZN(n51));
   AND2_X1 U53 (.A1(A[10]),
	.A2(n53),
	.ZN(n52));
   AND2_X1 U54 (.A1(A[9]),
	.A2(n54),
	.ZN(n53));
   AND2_X1 U55 (.A1(A[8]),
	.A2(n55),
	.ZN(n54));
   AND2_X1 U56 (.A1(A[7]),
	.A2(n30),
	.ZN(n55));
   AND2_X1 U57 (.A1(A[3]),
	.A2(A[2]),
	.ZN(n56));
   INV_X1 U58 (.A(A[2]),
	.ZN(SUM[2]));
endmodule

module fetch_unit (
	clk, 
	rst, 
	en, 
	PC_MUX_SEL, 
	IRAM_DOUT_IN, 
	PC_JUMP_ADDR, 
	PC, 
	IR_IN);
   input clk;
   input rst;
   input en;
   input PC_MUX_SEL;
   input [31:0] IRAM_DOUT_IN;
   input [31:0] PC_JUMP_ADDR;
   output [31:0] PC;
   output [31:0] IR_IN;

   // Internal wires
   wire FE_OFN37_n38;
   wire FE_OFN36_n37;
   wire N38;
   wire N39;
   wire N40;
   wire N41;
   wire N42;
   wire N43;
   wire N44;
   wire N45;
   wire N46;
   wire N47;
   wire N48;
   wire N49;
   wire N50;
   wire N51;
   wire N52;
   wire N53;
   wire N54;
   wire N55;
   wire N56;
   wire N57;
   wire N58;
   wire N59;
   wire N60;
   wire N61;
   wire N62;
   wire N63;
   wire N64;
   wire N65;
   wire N66;
   wire N67;
   wire N68;
   wire N69;
   wire n37;
   wire n38;
   wire n39;
   wire n41;
   wire n42;
   wire n43;
   wire n44;
   wire n45;
   wire n46;
   wire n47;
   wire n48;
   wire n49;
   wire n50;
   wire n51;
   wire n52;
   wire n53;
   wire n54;
   wire n55;
   wire n56;
   wire n57;
   wire n58;
   wire n59;
   wire n60;
   wire n61;
   wire n62;
   wire n63;
   wire n64;
   wire n65;
   wire n66;
   wire n67;
   wire n68;
   wire n69;
   wire n70;
   wire n71;
   wire n2;
   wire n3;
   wire n4;
   wire n5;
   wire n6;
   wire n7;
   wire n8;
   wire n9;
   wire n10;
   wire n20;
   wire n21;
   wire n22;
   wire n23;
   wire n24;
   wire n25;
   wire n26;
   wire n27;
   wire n28;
   wire n29;
   wire n30;
   wire n31;
   wire n32;
   wire n33;
   wire n34;
   wire n35;
   wire n36;
   wire n40;
   wire n72;
   wire n73;
   wire n74;
   wire n75;
   wire n76;
   wire n77;
   wire n78;
   wire n79;
   wire n80;
   wire n81;
   wire n82;
   wire n83;
   wire n84;

   assign IR_IN[31] = IRAM_DOUT_IN[31] ;
   assign IR_IN[30] = IRAM_DOUT_IN[30] ;
   assign IR_IN[29] = IRAM_DOUT_IN[29] ;
   assign IR_IN[28] = IRAM_DOUT_IN[28] ;
   assign IR_IN[27] = IRAM_DOUT_IN[27] ;
   assign IR_IN[26] = IRAM_DOUT_IN[26] ;
   assign IR_IN[25] = IRAM_DOUT_IN[25] ;
   assign IR_IN[24] = IRAM_DOUT_IN[24] ;
   assign IR_IN[23] = IRAM_DOUT_IN[23] ;
   assign IR_IN[22] = IRAM_DOUT_IN[22] ;
   assign IR_IN[21] = IRAM_DOUT_IN[21] ;
   assign IR_IN[20] = IRAM_DOUT_IN[20] ;
   assign IR_IN[19] = IRAM_DOUT_IN[19] ;
   assign IR_IN[18] = IRAM_DOUT_IN[18] ;
   assign IR_IN[17] = IRAM_DOUT_IN[17] ;
   assign IR_IN[16] = IRAM_DOUT_IN[16] ;
   assign IR_IN[15] = IRAM_DOUT_IN[15] ;
   assign IR_IN[14] = IRAM_DOUT_IN[14] ;
   assign IR_IN[13] = IRAM_DOUT_IN[13] ;
   assign IR_IN[12] = IRAM_DOUT_IN[12] ;
   assign IR_IN[11] = IRAM_DOUT_IN[11] ;
   assign IR_IN[10] = IRAM_DOUT_IN[10] ;
   assign IR_IN[9] = IRAM_DOUT_IN[9] ;
   assign IR_IN[8] = IRAM_DOUT_IN[8] ;
   assign IR_IN[7] = IRAM_DOUT_IN[7] ;
   assign IR_IN[6] = IRAM_DOUT_IN[6] ;
   assign IR_IN[5] = IRAM_DOUT_IN[5] ;
   assign IR_IN[4] = IRAM_DOUT_IN[4] ;
   assign IR_IN[3] = IRAM_DOUT_IN[3] ;
   assign IR_IN[2] = IRAM_DOUT_IN[2] ;
   assign IR_IN[1] = IRAM_DOUT_IN[1] ;
   assign IR_IN[0] = IRAM_DOUT_IN[0] ;

   BUF_X2 FE_OFC37_n38 (.A(n38),
	.Z(FE_OFN37_n38));
   BUF_X2 FE_OFC36_n37 (.A(n37),
	.Z(FE_OFN36_n37));
   DFF_X1 currPC_reg_0_ (.D(n83),
	.CK(clk),
	.Q(PC[0]));
   DFF_X1 currPC_reg_1_ (.D(n82),
	.CK(clk),
	.Q(PC[1]));
   DFF_X1 currPC_reg_2_ (.D(n81),
	.CK(clk),
	.Q(PC[2]));
   DFF_X1 currPC_reg_3_ (.D(n80),
	.CK(clk),
	.Q(PC[3]));
   DFF_X1 currPC_reg_4_ (.D(n79),
	.CK(clk),
	.Q(PC[4]));
   DFF_X1 currPC_reg_5_ (.D(n78),
	.CK(clk),
	.Q(PC[5]));
   DFF_X1 currPC_reg_6_ (.D(n77),
	.CK(clk),
	.Q(PC[6]));
   DFF_X1 currPC_reg_7_ (.D(n76),
	.CK(clk),
	.Q(PC[7]));
   DFF_X1 currPC_reg_8_ (.D(n75),
	.CK(clk),
	.Q(PC[8]));
   DFF_X1 currPC_reg_9_ (.D(n74),
	.CK(clk),
	.Q(PC[9]));
   DFF_X1 currPC_reg_10_ (.D(n73),
	.CK(clk),
	.Q(PC[10]));
   DFF_X1 currPC_reg_11_ (.D(n72),
	.CK(clk),
	.Q(PC[11]));
   DFF_X1 currPC_reg_12_ (.D(n40),
	.CK(clk),
	.Q(PC[12]));
   DFF_X1 currPC_reg_13_ (.D(n36),
	.CK(clk),
	.Q(PC[13]));
   DFF_X1 currPC_reg_14_ (.D(n35),
	.CK(clk),
	.Q(PC[14]));
   DFF_X1 currPC_reg_15_ (.D(n34),
	.CK(clk),
	.Q(PC[15]));
   DFF_X1 currPC_reg_16_ (.D(n33),
	.CK(clk),
	.Q(PC[16]));
   DFF_X1 currPC_reg_17_ (.D(n32),
	.CK(clk),
	.Q(PC[17]));
   DFF_X1 currPC_reg_18_ (.D(n31),
	.CK(clk),
	.Q(PC[18]));
   DFF_X1 currPC_reg_19_ (.D(n30),
	.CK(clk),
	.Q(PC[19]));
   DFF_X1 currPC_reg_20_ (.D(n29),
	.CK(clk),
	.Q(PC[20]));
   DFF_X1 currPC_reg_21_ (.D(n28),
	.CK(clk),
	.Q(PC[21]));
   DFF_X1 currPC_reg_22_ (.D(n27),
	.CK(clk),
	.Q(PC[22]));
   DFF_X1 currPC_reg_23_ (.D(n26),
	.CK(clk),
	.Q(PC[23]));
   DFF_X1 currPC_reg_24_ (.D(n25),
	.CK(clk),
	.Q(PC[24]));
   DFF_X1 currPC_reg_25_ (.D(n24),
	.CK(clk),
	.Q(PC[25]));
   DFF_X1 currPC_reg_26_ (.D(n23),
	.CK(clk),
	.Q(PC[26]));
   DFF_X1 currPC_reg_27_ (.D(n22),
	.CK(clk),
	.Q(PC[27]));
   DFF_X1 currPC_reg_28_ (.D(n21),
	.CK(clk),
	.Q(PC[28]));
   DFF_X1 currPC_reg_29_ (.D(n20),
	.CK(clk),
	.Q(PC[29]));
   DFF_X1 currPC_reg_30_ (.D(n3),
	.CK(clk),
	.Q(PC[30]));
   fetch_unit_DW01_add_0 add_33 (.A(PC),
	.B({ 1'b0,
		1'b0,
		1'b0,
		1'b0,
		1'b0,
		1'b0,
		1'b0,
		1'b0,
		1'b0,
		1'b0,
		1'b0,
		1'b0,
		1'b0,
		1'b0,
		1'b0,
		1'b0,
		1'b0,
		1'b0,
		1'b0,
		1'b0,
		1'b0,
		1'b0,
		1'b0,
		1'b0,
		1'b0,
		1'b0,
		1'b0,
		1'b0,
		1'b0,
		1'b1,
		1'b0,
		1'b0 }),
	.CI(1'b0),
	.SUM({ N69,
		N68,
		N67,
		N66,
		N65,
		N64,
		N63,
		N62,
		N61,
		N60,
		N59,
		N58,
		N57,
		N56,
		N55,
		N54,
		N53,
		N52,
		N51,
		N50,
		N49,
		N48,
		N47,
		N46,
		N45,
		N44,
		N43,
		N42,
		N41,
		N40,
		N39,
		N38 }));
   DFF_X1 currPC_reg_31_ (.D(n7),
	.CK(clk),
	.Q(PC[31]));
   AND2_X1 U4 (.A1(n9),
	.A2(n8),
	.ZN(n2));
   NAND3_X1 U6 (.A1(n4),
	.A2(n5),
	.A3(n6),
	.ZN(n3));
   NAND2_X1 U7 (.A1(n10),
	.A2(n2),
	.ZN(n7));
   NAND2_X1 U8 (.A1(PC[30]),
	.A2(FE_OFN36_n37),
	.ZN(n4));
   NAND2_X1 U9 (.A1(N68),
	.A2(FE_OFN37_n38),
	.ZN(n5));
   NAND2_X1 U10 (.A1(PC_JUMP_ADDR[30]),
	.A2(n39),
	.ZN(n6));
   NAND2_X1 U11 (.A1(PC[31]),
	.A2(FE_OFN36_n37),
	.ZN(n8));
   NAND2_X1 U12 (.A1(N69),
	.A2(FE_OFN37_n38),
	.ZN(n9));
   NAND2_X1 U13 (.A1(PC_JUMP_ADDR[31]),
	.A2(n39),
	.ZN(n10));
   NOR2_X1 U19 (.A1(n84),
	.A2(PC_MUX_SEL),
	.ZN(n38));
   INV_X1 U20 (.A(n71),
	.ZN(n84));
   AND2_X2 U22 (.A1(PC_MUX_SEL),
	.A2(n71),
	.ZN(n39));
   INV_X1 U25 (.A(n41),
	.ZN(n20));
   AOI222_X1 U26 (.A1(PC[29]),
	.A2(FE_OFN36_n37),
	.B1(N67),
	.B2(FE_OFN37_n38),
	.C1(PC_JUMP_ADDR[29]),
	.C2(n39),
	.ZN(n41));
   INV_X1 U27 (.A(n42),
	.ZN(n21));
   AOI222_X1 U28 (.A1(PC[28]),
	.A2(FE_OFN36_n37),
	.B1(N66),
	.B2(FE_OFN37_n38),
	.C1(PC_JUMP_ADDR[28]),
	.C2(n39),
	.ZN(n42));
   INV_X1 U29 (.A(n43),
	.ZN(n22));
   AOI222_X1 U30 (.A1(PC[27]),
	.A2(FE_OFN36_n37),
	.B1(N65),
	.B2(FE_OFN37_n38),
	.C1(PC_JUMP_ADDR[27]),
	.C2(n39),
	.ZN(n43));
   INV_X1 U31 (.A(n44),
	.ZN(n23));
   AOI222_X1 U32 (.A1(PC[26]),
	.A2(FE_OFN36_n37),
	.B1(N64),
	.B2(FE_OFN37_n38),
	.C1(PC_JUMP_ADDR[26]),
	.C2(n39),
	.ZN(n44));
   INV_X1 U33 (.A(n45),
	.ZN(n24));
   AOI222_X1 U34 (.A1(PC[25]),
	.A2(FE_OFN36_n37),
	.B1(N63),
	.B2(FE_OFN37_n38),
	.C1(PC_JUMP_ADDR[25]),
	.C2(n39),
	.ZN(n45));
   INV_X1 U35 (.A(n46),
	.ZN(n25));
   AOI222_X1 U36 (.A1(PC[24]),
	.A2(FE_OFN36_n37),
	.B1(N62),
	.B2(FE_OFN37_n38),
	.C1(PC_JUMP_ADDR[24]),
	.C2(n39),
	.ZN(n46));
   INV_X1 U37 (.A(n47),
	.ZN(n26));
   AOI222_X1 U38 (.A1(PC[23]),
	.A2(FE_OFN36_n37),
	.B1(N61),
	.B2(FE_OFN37_n38),
	.C1(PC_JUMP_ADDR[23]),
	.C2(n39),
	.ZN(n47));
   INV_X1 U39 (.A(n48),
	.ZN(n27));
   AOI222_X1 U40 (.A1(PC[22]),
	.A2(FE_OFN36_n37),
	.B1(N60),
	.B2(FE_OFN37_n38),
	.C1(PC_JUMP_ADDR[22]),
	.C2(n39),
	.ZN(n48));
   INV_X1 U41 (.A(n49),
	.ZN(n28));
   AOI222_X1 U42 (.A1(PC[21]),
	.A2(FE_OFN36_n37),
	.B1(N59),
	.B2(FE_OFN37_n38),
	.C1(PC_JUMP_ADDR[21]),
	.C2(n39),
	.ZN(n49));
   INV_X1 U43 (.A(n50),
	.ZN(n29));
   AOI222_X1 U44 (.A1(PC[20]),
	.A2(FE_OFN36_n37),
	.B1(N58),
	.B2(FE_OFN37_n38),
	.C1(PC_JUMP_ADDR[20]),
	.C2(n39),
	.ZN(n50));
   INV_X1 U45 (.A(n51),
	.ZN(n30));
   AOI222_X1 U46 (.A1(PC[19]),
	.A2(FE_OFN36_n37),
	.B1(N57),
	.B2(FE_OFN37_n38),
	.C1(PC_JUMP_ADDR[19]),
	.C2(n39),
	.ZN(n51));
   INV_X1 U47 (.A(n52),
	.ZN(n31));
   AOI222_X1 U48 (.A1(PC[18]),
	.A2(FE_OFN36_n37),
	.B1(N56),
	.B2(FE_OFN37_n38),
	.C1(PC_JUMP_ADDR[18]),
	.C2(n39),
	.ZN(n52));
   INV_X1 U49 (.A(n53),
	.ZN(n32));
   AOI222_X1 U50 (.A1(PC[17]),
	.A2(FE_OFN36_n37),
	.B1(N55),
	.B2(FE_OFN37_n38),
	.C1(PC_JUMP_ADDR[17]),
	.C2(n39),
	.ZN(n53));
   INV_X1 U51 (.A(n54),
	.ZN(n33));
   AOI222_X1 U52 (.A1(PC[16]),
	.A2(FE_OFN36_n37),
	.B1(N54),
	.B2(FE_OFN37_n38),
	.C1(PC_JUMP_ADDR[16]),
	.C2(n39),
	.ZN(n54));
   INV_X1 U53 (.A(n55),
	.ZN(n34));
   AOI222_X1 U54 (.A1(PC[15]),
	.A2(FE_OFN36_n37),
	.B1(N53),
	.B2(FE_OFN37_n38),
	.C1(PC_JUMP_ADDR[15]),
	.C2(n39),
	.ZN(n55));
   INV_X1 U55 (.A(n56),
	.ZN(n35));
   AOI222_X1 U56 (.A1(PC[14]),
	.A2(FE_OFN36_n37),
	.B1(N52),
	.B2(FE_OFN37_n38),
	.C1(PC_JUMP_ADDR[14]),
	.C2(n39),
	.ZN(n56));
   INV_X1 U57 (.A(n57),
	.ZN(n36));
   AOI222_X1 U58 (.A1(PC[13]),
	.A2(FE_OFN36_n37),
	.B1(N51),
	.B2(FE_OFN37_n38),
	.C1(PC_JUMP_ADDR[13]),
	.C2(n39),
	.ZN(n57));
   NOR2_X1 U59 (.A1(en),
	.A2(rst),
	.ZN(n37));
   NOR2_X1 U60 (.A1(FE_OFN36_n37),
	.A2(rst),
	.ZN(n71));
   INV_X1 U61 (.A(n58),
	.ZN(n40));
   AOI222_X1 U62 (.A1(PC[12]),
	.A2(FE_OFN36_n37),
	.B1(N50),
	.B2(FE_OFN37_n38),
	.C1(PC_JUMP_ADDR[12]),
	.C2(n39),
	.ZN(n58));
   INV_X1 U63 (.A(n59),
	.ZN(n72));
   AOI222_X1 U64 (.A1(PC[11]),
	.A2(FE_OFN36_n37),
	.B1(N49),
	.B2(FE_OFN37_n38),
	.C1(PC_JUMP_ADDR[11]),
	.C2(n39),
	.ZN(n59));
   INV_X1 U65 (.A(n60),
	.ZN(n73));
   AOI222_X1 U66 (.A1(PC[10]),
	.A2(FE_OFN36_n37),
	.B1(N48),
	.B2(FE_OFN37_n38),
	.C1(PC_JUMP_ADDR[10]),
	.C2(n39),
	.ZN(n60));
   INV_X1 U67 (.A(n61),
	.ZN(n74));
   AOI222_X1 U68 (.A1(PC[9]),
	.A2(FE_OFN36_n37),
	.B1(N47),
	.B2(FE_OFN37_n38),
	.C1(PC_JUMP_ADDR[9]),
	.C2(n39),
	.ZN(n61));
   INV_X1 U69 (.A(n62),
	.ZN(n75));
   AOI222_X1 U70 (.A1(PC[8]),
	.A2(FE_OFN36_n37),
	.B1(N46),
	.B2(FE_OFN37_n38),
	.C1(PC_JUMP_ADDR[8]),
	.C2(n39),
	.ZN(n62));
   INV_X1 U71 (.A(n63),
	.ZN(n76));
   AOI222_X1 U72 (.A1(PC[7]),
	.A2(FE_OFN36_n37),
	.B1(N45),
	.B2(FE_OFN37_n38),
	.C1(PC_JUMP_ADDR[7]),
	.C2(n39),
	.ZN(n63));
   INV_X1 U73 (.A(n64),
	.ZN(n77));
   AOI222_X1 U74 (.A1(PC[6]),
	.A2(FE_OFN36_n37),
	.B1(N44),
	.B2(FE_OFN37_n38),
	.C1(PC_JUMP_ADDR[6]),
	.C2(n39),
	.ZN(n64));
   INV_X1 U75 (.A(n65),
	.ZN(n78));
   AOI222_X1 U76 (.A1(PC[5]),
	.A2(FE_OFN36_n37),
	.B1(N43),
	.B2(FE_OFN37_n38),
	.C1(PC_JUMP_ADDR[5]),
	.C2(n39),
	.ZN(n65));
   INV_X1 U77 (.A(n66),
	.ZN(n79));
   AOI222_X1 U78 (.A1(PC[4]),
	.A2(FE_OFN36_n37),
	.B1(N42),
	.B2(FE_OFN37_n38),
	.C1(PC_JUMP_ADDR[4]),
	.C2(n39),
	.ZN(n66));
   INV_X1 U79 (.A(n67),
	.ZN(n80));
   AOI222_X1 U80 (.A1(PC[3]),
	.A2(FE_OFN36_n37),
	.B1(N41),
	.B2(FE_OFN37_n38),
	.C1(PC_JUMP_ADDR[3]),
	.C2(n39),
	.ZN(n67));
   INV_X1 U81 (.A(n68),
	.ZN(n81));
   AOI222_X1 U82 (.A1(PC[2]),
	.A2(FE_OFN36_n37),
	.B1(N40),
	.B2(FE_OFN37_n38),
	.C1(PC_JUMP_ADDR[2]),
	.C2(n39),
	.ZN(n68));
   INV_X1 U83 (.A(n69),
	.ZN(n82));
   AOI222_X1 U84 (.A1(PC[1]),
	.A2(FE_OFN36_n37),
	.B1(N39),
	.B2(FE_OFN37_n38),
	.C1(PC_JUMP_ADDR[1]),
	.C2(n39),
	.ZN(n69));
   INV_X1 U85 (.A(n70),
	.ZN(n83));
   AOI222_X1 U86 (.A1(PC[0]),
	.A2(FE_OFN36_n37),
	.B1(N38),
	.B2(FE_OFN37_n38),
	.C1(PC_JUMP_ADDR[0]),
	.C2(n39),
	.ZN(n70));
endmodule

module register_file_NBITS32 (
	CLK, 
	RESET, 
	ENABLE, 
	RD1, 
	RD2, 
	WR, 
	ADD_WR, 
	ADD_RD1, 
	ADD_RD2, 
	DATAIN, 
	OUT1, 
	OUT2);
   input CLK;
   input RESET;
   input ENABLE;
   input RD1;
   input RD2;
   input WR;
   input [4:0] ADD_WR;
   input [4:0] ADD_RD1;
   input [4:0] ADD_RD2;
   input [31:0] DATAIN;
   output [31:0] OUT1;
   output [31:0] OUT2;

   // Internal wires
   wire FE_OFN136_n2761;
   wire FE_OFN135_n2761;
   wire FE_OFN134_n3573;
   wire FE_OFN133_n3573;
   wire FE_OFN132_n3570;
   wire FE_OFN131_n3570;
   wire FE_OFN114_n2768;
   wire FE_OFN113_n2768;
   wire FE_OFN112_n2763;
   wire FE_OFN111_n2763;
   wire FE_OFN110_n2763;
   wire FE_OFN109_n3569;
   wire FE_OFN108_n3569;
   wire FE_OFN107_n3576;
   wire FE_OFN106_n3576;
   wire FE_OFN105_n3576;
   wire FE_OFN89_n4027;
   wire FE_OFN88_n4010;
   wire FE_OFN87_n4032;
   wire FE_OFN86_n4008;
   wire FE_OFN85_n4022;
   wire FE_OFN84_n4005;
   wire FE_OFN83_n4024;
   wire FE_OFN82_n4007;
   wire FE_OFN81_n4030;
   wire FE_OFN80_n4035;
   wire FE_OFN79_n4023;
   wire FE_OFN78_n4014;
   wire FE_OFN77_n4026;
   wire FE_OFN76_n4013;
   wire FE_OFN75_n4028;
   wire FE_OFN74_n4015;
   wire FE_OFN73_n4009;
   wire FE_OFN72_n4021;
   wire FE_OFN71_n4006;
   wire FE_OFN70_n4033;
   wire FE_OFN69_n4025;
   wire FE_OFN68_n4011;
   wire FE_OFN67_n4029;
   wire FE_OFN66_n4017;
   wire FE_OFN65_n4018;
   wire FE_OFN64_n4012;
   wire FE_OFN63_n4031;
   wire FE_OFN62_n4016;
   wire FE_OFN61_n4019;
   wire FE_OFN60_n4036;
   wire FE_OFN59_n4034;
   wire FE_OFN56_n2764;
   wire FE_OFN55_n2764;
   wire FE_OFN54_n2764;
   wire FE_OFN53_n2765;
   wire FE_OFN52_n2765;
   wire FE_OFN51_n2765;
   wire FE_OFN50_n3575;
   wire FE_OFN49_n3575;
   wire FE_OFN48_n3575;
   wire FE_OFN47_n3572;
   wire FE_OFN46_n3572;
   wire FE_OFN38_n3588;
   wire FE_OFN33_n3584;
   wire FE_OFN32_n2776;
   wire FE_OFN31_n3582;
   wire FE_OFN30_n2774;
   wire FE_OFN18_n4041;
   wire FE_OFN14_n2762;
   wire FE_OFN13_n2762;
   wire FE_OFN12_n2767;
   wire FE_OFN11_n2767;
   wire FE_OFN10_n2766;
   wire FE_OFN9_n2766;
   wire FE_OFN8_n2766;
   wire FE_OFN7_n3571;
   wire FE_OFN6_n3571;
   wire FE_OFN5_n3574;
   wire FE_OFN4_n3574;
   wire FE_OFN3_n3574;
   wire N31;
   wire N32;
   wire N33;
   wire N34;
   wire N35;
   wire N36;
   wire N37;
   wire N38;
   wire N39;
   wire N40;
   wire N41;
   wire N42;
   wire N43;
   wire N44;
   wire N45;
   wire N46;
   wire N47;
   wire N48;
   wire N49;
   wire N50;
   wire N51;
   wire N52;
   wire N53;
   wire N54;
   wire N55;
   wire N56;
   wire N57;
   wire N58;
   wire N59;
   wire N60;
   wire N61;
   wire N62;
   wire N96;
   wire N97;
   wire N98;
   wire N99;
   wire N100;
   wire N101;
   wire N102;
   wire N103;
   wire N104;
   wire N105;
   wire N106;
   wire N107;
   wire N108;
   wire N109;
   wire N110;
   wire N111;
   wire N112;
   wire N113;
   wire N114;
   wire N115;
   wire N116;
   wire N117;
   wire N118;
   wire N119;
   wire N120;
   wire N121;
   wire N122;
   wire N123;
   wire N124;
   wire N125;
   wire N126;
   wire N127;
   wire n38;
   wire n39;
   wire n40;
   wire n41;
   wire n42;
   wire n43;
   wire n44;
   wire n45;
   wire n46;
   wire n47;
   wire n48;
   wire n49;
   wire n50;
   wire n51;
   wire n52;
   wire n53;
   wire n54;
   wire n55;
   wire n56;
   wire n57;
   wire n58;
   wire n59;
   wire n60;
   wire n61;
   wire n62;
   wire n63;
   wire n64;
   wire n65;
   wire n66;
   wire n67;
   wire n68;
   wire n69;
   wire n70;
   wire n71;
   wire n72;
   wire n73;
   wire n74;
   wire n75;
   wire n76;
   wire n77;
   wire n78;
   wire n79;
   wire n80;
   wire n81;
   wire n82;
   wire n83;
   wire n84;
   wire n85;
   wire n86;
   wire n87;
   wire n88;
   wire n89;
   wire n90;
   wire n91;
   wire n92;
   wire n93;
   wire n94;
   wire n95;
   wire n96;
   wire n97;
   wire n98;
   wire n99;
   wire n100;
   wire n101;
   wire n102;
   wire n103;
   wire n104;
   wire n105;
   wire n106;
   wire n107;
   wire n108;
   wire n109;
   wire n110;
   wire n111;
   wire n112;
   wire n113;
   wire n114;
   wire n115;
   wire n116;
   wire n117;
   wire n118;
   wire n119;
   wire n120;
   wire n121;
   wire n122;
   wire n123;
   wire n124;
   wire n125;
   wire n126;
   wire n127;
   wire n128;
   wire n129;
   wire n130;
   wire n131;
   wire n132;
   wire n133;
   wire n134;
   wire n135;
   wire n136;
   wire n137;
   wire n138;
   wire n139;
   wire n140;
   wire n141;
   wire n142;
   wire n143;
   wire n144;
   wire n145;
   wire n146;
   wire n147;
   wire n148;
   wire n149;
   wire n150;
   wire n151;
   wire n152;
   wire n153;
   wire n154;
   wire n155;
   wire n156;
   wire n157;
   wire n158;
   wire n159;
   wire n160;
   wire n161;
   wire n162;
   wire n163;
   wire n164;
   wire n165;
   wire n166;
   wire n167;
   wire n168;
   wire n169;
   wire n170;
   wire n171;
   wire n172;
   wire n173;
   wire n174;
   wire n175;
   wire n176;
   wire n177;
   wire n178;
   wire n179;
   wire n180;
   wire n181;
   wire n182;
   wire n183;
   wire n184;
   wire n185;
   wire n186;
   wire n187;
   wire n188;
   wire n189;
   wire n190;
   wire n191;
   wire n192;
   wire n193;
   wire n194;
   wire n195;
   wire n196;
   wire n197;
   wire n198;
   wire n199;
   wire n200;
   wire n201;
   wire n202;
   wire n203;
   wire n204;
   wire n205;
   wire n206;
   wire n207;
   wire n208;
   wire n209;
   wire n210;
   wire n211;
   wire n212;
   wire n213;
   wire n214;
   wire n215;
   wire n216;
   wire n217;
   wire n218;
   wire n219;
   wire n220;
   wire n221;
   wire n222;
   wire n223;
   wire n224;
   wire n225;
   wire n226;
   wire n227;
   wire n228;
   wire n229;
   wire n230;
   wire n231;
   wire n232;
   wire n233;
   wire n234;
   wire n235;
   wire n236;
   wire n237;
   wire n238;
   wire n239;
   wire n240;
   wire n241;
   wire n242;
   wire n243;
   wire n244;
   wire n245;
   wire n246;
   wire n247;
   wire n248;
   wire n249;
   wire n250;
   wire n251;
   wire n252;
   wire n253;
   wire n254;
   wire n255;
   wire n256;
   wire n257;
   wire n258;
   wire n259;
   wire n260;
   wire n261;
   wire n262;
   wire n263;
   wire n264;
   wire n265;
   wire n266;
   wire n267;
   wire n268;
   wire n269;
   wire n270;
   wire n271;
   wire n272;
   wire n273;
   wire n274;
   wire n275;
   wire n276;
   wire n277;
   wire n278;
   wire n279;
   wire n280;
   wire n281;
   wire n282;
   wire n283;
   wire n284;
   wire n285;
   wire n286;
   wire n287;
   wire n288;
   wire n289;
   wire n290;
   wire n291;
   wire n292;
   wire n293;
   wire n294;
   wire n295;
   wire n296;
   wire n297;
   wire n298;
   wire n299;
   wire n300;
   wire n301;
   wire n302;
   wire n303;
   wire n304;
   wire n305;
   wire n306;
   wire n307;
   wire n308;
   wire n309;
   wire n310;
   wire n311;
   wire n312;
   wire n313;
   wire n314;
   wire n315;
   wire n316;
   wire n317;
   wire n318;
   wire n319;
   wire n320;
   wire n321;
   wire n322;
   wire n323;
   wire n324;
   wire n325;
   wire n326;
   wire n327;
   wire n328;
   wire n329;
   wire n330;
   wire n331;
   wire n332;
   wire n333;
   wire n334;
   wire n335;
   wire n336;
   wire n337;
   wire n338;
   wire n339;
   wire n340;
   wire n341;
   wire n342;
   wire n343;
   wire n344;
   wire n345;
   wire n346;
   wire n347;
   wire n348;
   wire n349;
   wire n350;
   wire n351;
   wire n352;
   wire n353;
   wire n354;
   wire n355;
   wire n356;
   wire n357;
   wire n358;
   wire n359;
   wire n360;
   wire n361;
   wire n362;
   wire n363;
   wire n364;
   wire n365;
   wire n366;
   wire n367;
   wire n368;
   wire n369;
   wire n370;
   wire n371;
   wire n372;
   wire n373;
   wire n374;
   wire n375;
   wire n376;
   wire n377;
   wire n378;
   wire n379;
   wire n380;
   wire n381;
   wire n382;
   wire n383;
   wire n384;
   wire n385;
   wire n386;
   wire n387;
   wire n388;
   wire n389;
   wire n390;
   wire n391;
   wire n392;
   wire n393;
   wire n394;
   wire n395;
   wire n396;
   wire n397;
   wire n398;
   wire n399;
   wire n400;
   wire n401;
   wire n402;
   wire n403;
   wire n404;
   wire n405;
   wire n406;
   wire n407;
   wire n408;
   wire n409;
   wire n410;
   wire n411;
   wire n412;
   wire n413;
   wire n414;
   wire n415;
   wire n416;
   wire n417;
   wire n418;
   wire n419;
   wire n420;
   wire n421;
   wire n422;
   wire n423;
   wire n424;
   wire n425;
   wire n426;
   wire n427;
   wire n428;
   wire n429;
   wire n430;
   wire n431;
   wire n432;
   wire n433;
   wire n434;
   wire n435;
   wire n436;
   wire n437;
   wire n438;
   wire n439;
   wire n440;
   wire n441;
   wire n442;
   wire n443;
   wire n444;
   wire n445;
   wire n446;
   wire n447;
   wire n448;
   wire n449;
   wire n450;
   wire n451;
   wire n452;
   wire n453;
   wire n454;
   wire n455;
   wire n456;
   wire n457;
   wire n458;
   wire n459;
   wire n460;
   wire n461;
   wire n462;
   wire n463;
   wire n464;
   wire n465;
   wire n466;
   wire n467;
   wire n468;
   wire n469;
   wire n470;
   wire n471;
   wire n472;
   wire n473;
   wire n474;
   wire n475;
   wire n476;
   wire n477;
   wire n478;
   wire n479;
   wire n480;
   wire n481;
   wire n482;
   wire n483;
   wire n484;
   wire n485;
   wire n486;
   wire n487;
   wire n488;
   wire n489;
   wire n490;
   wire n491;
   wire n492;
   wire n493;
   wire n494;
   wire n495;
   wire n496;
   wire n497;
   wire n498;
   wire n499;
   wire n500;
   wire n501;
   wire n502;
   wire n503;
   wire n504;
   wire n505;
   wire n506;
   wire n507;
   wire n508;
   wire n509;
   wire n510;
   wire n511;
   wire n512;
   wire n513;
   wire n514;
   wire n515;
   wire n516;
   wire n517;
   wire n518;
   wire n519;
   wire n520;
   wire n521;
   wire n522;
   wire n523;
   wire n524;
   wire n525;
   wire n526;
   wire n527;
   wire n528;
   wire n529;
   wire n530;
   wire n531;
   wire n532;
   wire n533;
   wire n534;
   wire n535;
   wire n536;
   wire n537;
   wire n538;
   wire n539;
   wire n540;
   wire n541;
   wire n542;
   wire n543;
   wire n544;
   wire n545;
   wire n546;
   wire n547;
   wire n548;
   wire n549;
   wire n550;
   wire n551;
   wire n552;
   wire n553;
   wire n554;
   wire n555;
   wire n556;
   wire n557;
   wire n558;
   wire n559;
   wire n560;
   wire n561;
   wire n562;
   wire n563;
   wire n564;
   wire n565;
   wire n566;
   wire n567;
   wire n568;
   wire n569;
   wire n570;
   wire n571;
   wire n572;
   wire n573;
   wire n574;
   wire n575;
   wire n576;
   wire n577;
   wire n578;
   wire n579;
   wire n580;
   wire n581;
   wire n582;
   wire n583;
   wire n584;
   wire n585;
   wire n586;
   wire n587;
   wire n588;
   wire n589;
   wire n590;
   wire n591;
   wire n592;
   wire n593;
   wire n594;
   wire n595;
   wire n596;
   wire n597;
   wire n598;
   wire n599;
   wire n600;
   wire n601;
   wire n602;
   wire n603;
   wire n604;
   wire n605;
   wire n606;
   wire n607;
   wire n608;
   wire n609;
   wire n610;
   wire n611;
   wire n612;
   wire n613;
   wire n614;
   wire n615;
   wire n616;
   wire n617;
   wire n618;
   wire n619;
   wire n620;
   wire n621;
   wire n622;
   wire n623;
   wire n624;
   wire n625;
   wire n626;
   wire n627;
   wire n628;
   wire n629;
   wire n630;
   wire n631;
   wire n632;
   wire n633;
   wire n634;
   wire n635;
   wire n636;
   wire n637;
   wire n638;
   wire n639;
   wire n640;
   wire n641;
   wire n642;
   wire n643;
   wire n644;
   wire n645;
   wire n646;
   wire n647;
   wire n648;
   wire n649;
   wire n650;
   wire n651;
   wire n652;
   wire n653;
   wire n654;
   wire n655;
   wire n656;
   wire n657;
   wire n658;
   wire n659;
   wire n660;
   wire n661;
   wire n662;
   wire n663;
   wire n664;
   wire n665;
   wire n666;
   wire n667;
   wire n668;
   wire n669;
   wire n670;
   wire n671;
   wire n672;
   wire n673;
   wire n674;
   wire n675;
   wire n676;
   wire n677;
   wire n678;
   wire n679;
   wire n680;
   wire n681;
   wire n682;
   wire n683;
   wire n684;
   wire n685;
   wire n686;
   wire n687;
   wire n688;
   wire n689;
   wire n690;
   wire n691;
   wire n692;
   wire n693;
   wire n694;
   wire n695;
   wire n696;
   wire n697;
   wire n698;
   wire n699;
   wire n700;
   wire n701;
   wire n702;
   wire n703;
   wire n704;
   wire n705;
   wire n706;
   wire n707;
   wire n708;
   wire n709;
   wire n710;
   wire n711;
   wire n712;
   wire n713;
   wire n714;
   wire n715;
   wire n716;
   wire n717;
   wire n718;
   wire n719;
   wire n720;
   wire n721;
   wire n722;
   wire n723;
   wire n724;
   wire n725;
   wire n726;
   wire n727;
   wire n728;
   wire n729;
   wire n730;
   wire n731;
   wire n732;
   wire n733;
   wire n734;
   wire n735;
   wire n736;
   wire n737;
   wire n738;
   wire n739;
   wire n740;
   wire n741;
   wire n742;
   wire n743;
   wire n744;
   wire n745;
   wire n746;
   wire n747;
   wire n748;
   wire n749;
   wire n750;
   wire n751;
   wire n752;
   wire n753;
   wire n754;
   wire n755;
   wire n756;
   wire n757;
   wire n758;
   wire n759;
   wire n760;
   wire n761;
   wire n762;
   wire n763;
   wire n764;
   wire n765;
   wire n766;
   wire n767;
   wire n768;
   wire n769;
   wire n770;
   wire n771;
   wire n772;
   wire n773;
   wire n774;
   wire n775;
   wire n776;
   wire n777;
   wire n778;
   wire n779;
   wire n780;
   wire n781;
   wire n782;
   wire n783;
   wire n784;
   wire n785;
   wire n786;
   wire n787;
   wire n788;
   wire n789;
   wire n790;
   wire n791;
   wire n792;
   wire n793;
   wire n794;
   wire n795;
   wire n796;
   wire n797;
   wire n798;
   wire n799;
   wire n800;
   wire n801;
   wire n802;
   wire n803;
   wire n804;
   wire n805;
   wire n806;
   wire n807;
   wire n808;
   wire n809;
   wire n810;
   wire n811;
   wire n812;
   wire n813;
   wire n814;
   wire n815;
   wire n816;
   wire n817;
   wire n818;
   wire n819;
   wire n820;
   wire n821;
   wire n822;
   wire n823;
   wire n824;
   wire n825;
   wire n826;
   wire n827;
   wire n828;
   wire n829;
   wire n830;
   wire n831;
   wire n832;
   wire n833;
   wire n834;
   wire n835;
   wire n836;
   wire n837;
   wire n838;
   wire n839;
   wire n840;
   wire n841;
   wire n842;
   wire n843;
   wire n844;
   wire n845;
   wire n846;
   wire n847;
   wire n848;
   wire n849;
   wire n850;
   wire n851;
   wire n852;
   wire n853;
   wire n854;
   wire n855;
   wire n856;
   wire n857;
   wire n858;
   wire n859;
   wire n860;
   wire n861;
   wire n862;
   wire n863;
   wire n864;
   wire n865;
   wire n866;
   wire n867;
   wire n868;
   wire n869;
   wire n870;
   wire n871;
   wire n872;
   wire n873;
   wire n874;
   wire n875;
   wire n876;
   wire n877;
   wire n878;
   wire n879;
   wire n880;
   wire n881;
   wire n882;
   wire n883;
   wire n884;
   wire n885;
   wire n886;
   wire n887;
   wire n888;
   wire n889;
   wire n890;
   wire n891;
   wire n892;
   wire n893;
   wire n894;
   wire n895;
   wire n896;
   wire n897;
   wire n898;
   wire n899;
   wire n900;
   wire n901;
   wire n902;
   wire n903;
   wire n904;
   wire n905;
   wire n906;
   wire n907;
   wire n908;
   wire n909;
   wire n910;
   wire n911;
   wire n912;
   wire n913;
   wire n914;
   wire n915;
   wire n916;
   wire n917;
   wire n918;
   wire n919;
   wire n920;
   wire n921;
   wire n922;
   wire n923;
   wire n924;
   wire n925;
   wire n926;
   wire n927;
   wire n928;
   wire n929;
   wire n930;
   wire n931;
   wire n932;
   wire n933;
   wire n934;
   wire n935;
   wire n936;
   wire n937;
   wire n938;
   wire n939;
   wire n940;
   wire n941;
   wire n942;
   wire n943;
   wire n944;
   wire n945;
   wire n946;
   wire n947;
   wire n948;
   wire n949;
   wire n950;
   wire n951;
   wire n952;
   wire n953;
   wire n954;
   wire n955;
   wire n956;
   wire n957;
   wire n958;
   wire n959;
   wire n960;
   wire n961;
   wire n962;
   wire n963;
   wire n964;
   wire n965;
   wire n966;
   wire n967;
   wire n968;
   wire n969;
   wire n970;
   wire n971;
   wire n972;
   wire n973;
   wire n974;
   wire n975;
   wire n976;
   wire n977;
   wire n978;
   wire n979;
   wire n980;
   wire n981;
   wire n982;
   wire n983;
   wire n984;
   wire n985;
   wire n986;
   wire n987;
   wire n988;
   wire n989;
   wire n990;
   wire n991;
   wire n992;
   wire n993;
   wire n994;
   wire n995;
   wire n996;
   wire n997;
   wire n998;
   wire n999;
   wire n1000;
   wire n1001;
   wire n1002;
   wire n1003;
   wire n1004;
   wire n1005;
   wire n1006;
   wire n1007;
   wire n1008;
   wire n1009;
   wire n1010;
   wire n1011;
   wire n1012;
   wire n1013;
   wire n1014;
   wire n1015;
   wire n1016;
   wire n1017;
   wire n1018;
   wire n1019;
   wire n1020;
   wire n1021;
   wire n1022;
   wire n1023;
   wire n1024;
   wire n1025;
   wire n1026;
   wire n1027;
   wire n1028;
   wire n1029;
   wire n1030;
   wire n1031;
   wire n1032;
   wire n1033;
   wire n1034;
   wire n1035;
   wire n1036;
   wire n1037;
   wire n1038;
   wire n1039;
   wire n1040;
   wire n1041;
   wire n1042;
   wire n1043;
   wire n1044;
   wire n1045;
   wire n1046;
   wire n1047;
   wire n1048;
   wire n1049;
   wire n1050;
   wire n1051;
   wire n1052;
   wire n1053;
   wire n1054;
   wire n1055;
   wire n1056;
   wire n1057;
   wire n1058;
   wire n1059;
   wire n1060;
   wire n1061;
   wire n1062;
   wire n1063;
   wire n1064;
   wire n1065;
   wire n1066;
   wire n1067;
   wire n1068;
   wire n1069;
   wire n1070;
   wire n1071;
   wire n1072;
   wire n1073;
   wire n1074;
   wire n1075;
   wire n1076;
   wire n1077;
   wire n1078;
   wire n1079;
   wire n1080;
   wire n1081;
   wire n1082;
   wire n1083;
   wire n1084;
   wire n1085;
   wire n1086;
   wire n1087;
   wire n1088;
   wire n1089;
   wire n1090;
   wire n1091;
   wire n1092;
   wire n1093;
   wire n1094;
   wire n1095;
   wire n1096;
   wire n1097;
   wire n1098;
   wire n1099;
   wire n1100;
   wire n1101;
   wire n1102;
   wire n1103;
   wire n1104;
   wire n1105;
   wire n1106;
   wire n1107;
   wire n1108;
   wire n1109;
   wire n1110;
   wire n1111;
   wire n1112;
   wire n1113;
   wire n1114;
   wire n1115;
   wire n1116;
   wire n1117;
   wire n1118;
   wire n1119;
   wire n1120;
   wire n1121;
   wire n1122;
   wire n1123;
   wire n1124;
   wire n1125;
   wire n1126;
   wire n1127;
   wire n1128;
   wire n1129;
   wire n1130;
   wire n1131;
   wire n1132;
   wire n1133;
   wire n1134;
   wire n1135;
   wire n1136;
   wire n1137;
   wire n1138;
   wire n1139;
   wire n1140;
   wire n1141;
   wire n1142;
   wire n1143;
   wire n1144;
   wire n1145;
   wire n1146;
   wire n1147;
   wire n1148;
   wire n1149;
   wire n1150;
   wire n1151;
   wire n1152;
   wire n1153;
   wire n1154;
   wire n1155;
   wire n1156;
   wire n1157;
   wire n1158;
   wire n1159;
   wire n1160;
   wire n1161;
   wire n1162;
   wire n1163;
   wire n1164;
   wire n1165;
   wire n1166;
   wire n1167;
   wire n1168;
   wire n1169;
   wire n1170;
   wire n1171;
   wire n1172;
   wire n1173;
   wire n1174;
   wire n1175;
   wire n1176;
   wire n1177;
   wire n1178;
   wire n1179;
   wire n1180;
   wire n1181;
   wire n1182;
   wire n1183;
   wire n1184;
   wire n1185;
   wire n1186;
   wire n1187;
   wire n1188;
   wire n1189;
   wire n1190;
   wire n1191;
   wire n1192;
   wire n1193;
   wire n1194;
   wire n1195;
   wire n1196;
   wire n1197;
   wire n1198;
   wire n1199;
   wire n1200;
   wire n1201;
   wire n1202;
   wire n1203;
   wire n1204;
   wire n1205;
   wire n1206;
   wire n1207;
   wire n1208;
   wire n1209;
   wire n1210;
   wire n1211;
   wire n1212;
   wire n1213;
   wire n1214;
   wire n1215;
   wire n1216;
   wire n1217;
   wire n1218;
   wire n1219;
   wire n1220;
   wire n1221;
   wire n1222;
   wire n1223;
   wire n1224;
   wire n1225;
   wire n1226;
   wire n1227;
   wire n1228;
   wire n1229;
   wire n1230;
   wire n1231;
   wire n1232;
   wire n1233;
   wire n1234;
   wire n1235;
   wire n1236;
   wire n1237;
   wire n1238;
   wire n1239;
   wire n1240;
   wire n1241;
   wire n1242;
   wire n1243;
   wire n1244;
   wire n1245;
   wire n1246;
   wire n1247;
   wire n1248;
   wire n1249;
   wire n1250;
   wire n1251;
   wire n1252;
   wire n1253;
   wire n1254;
   wire n1255;
   wire n1256;
   wire n1257;
   wire n1258;
   wire n1259;
   wire n1260;
   wire n1261;
   wire n1262;
   wire n1263;
   wire n1264;
   wire n1265;
   wire n1266;
   wire n1267;
   wire n1268;
   wire n1269;
   wire n1270;
   wire n1271;
   wire n1272;
   wire n1273;
   wire n1274;
   wire n1275;
   wire n1276;
   wire n1277;
   wire n1278;
   wire n1279;
   wire n1280;
   wire n1281;
   wire n1282;
   wire n1283;
   wire n1284;
   wire n1285;
   wire n1286;
   wire n1287;
   wire n1288;
   wire n1289;
   wire n1290;
   wire n1291;
   wire n1292;
   wire n1293;
   wire n1294;
   wire n1295;
   wire n1296;
   wire n1297;
   wire n1298;
   wire n1299;
   wire n1300;
   wire n1301;
   wire n1302;
   wire n1303;
   wire n1304;
   wire n1305;
   wire n1306;
   wire n1307;
   wire n1308;
   wire n1309;
   wire n1310;
   wire n1311;
   wire n1312;
   wire n1313;
   wire n1314;
   wire n1315;
   wire n1316;
   wire n1317;
   wire n1318;
   wire n1319;
   wire n1320;
   wire n1321;
   wire n1322;
   wire n1323;
   wire n1324;
   wire n1325;
   wire n1326;
   wire n1327;
   wire n1328;
   wire n1329;
   wire n1330;
   wire n1331;
   wire n1332;
   wire n1333;
   wire n1334;
   wire n1335;
   wire n1336;
   wire n1337;
   wire n1338;
   wire n1339;
   wire n1340;
   wire n1341;
   wire n1342;
   wire n1343;
   wire n1344;
   wire n1345;
   wire n1346;
   wire n1347;
   wire n1348;
   wire n1349;
   wire n1350;
   wire n1351;
   wire n1352;
   wire n1353;
   wire n1354;
   wire n1355;
   wire n1356;
   wire n1357;
   wire n1358;
   wire n1359;
   wire n1360;
   wire n1361;
   wire n1362;
   wire n1363;
   wire n1364;
   wire n1365;
   wire n1366;
   wire n1367;
   wire n1368;
   wire n1369;
   wire n1370;
   wire n1371;
   wire n1372;
   wire n1373;
   wire n1374;
   wire n1375;
   wire n1376;
   wire n1377;
   wire n1378;
   wire n1379;
   wire n1380;
   wire n1381;
   wire n1382;
   wire n1383;
   wire n1384;
   wire n1385;
   wire n1386;
   wire n1387;
   wire n1388;
   wire n1389;
   wire n1390;
   wire n1391;
   wire n1392;
   wire n1393;
   wire n1394;
   wire n1395;
   wire n1396;
   wire n1397;
   wire n1398;
   wire n1399;
   wire n1400;
   wire n1401;
   wire n1402;
   wire n1403;
   wire n1404;
   wire n1405;
   wire n1406;
   wire n1407;
   wire n1408;
   wire n1409;
   wire n1410;
   wire n1411;
   wire n1412;
   wire n1413;
   wire n1414;
   wire n1415;
   wire n1416;
   wire n1417;
   wire n1418;
   wire n1419;
   wire n1420;
   wire n1421;
   wire n1422;
   wire n1423;
   wire n1424;
   wire n1425;
   wire n1426;
   wire n1427;
   wire n1428;
   wire n1429;
   wire n1430;
   wire n1431;
   wire n1432;
   wire n1433;
   wire n1434;
   wire n1435;
   wire n1436;
   wire n1437;
   wire n1438;
   wire n1439;
   wire n1440;
   wire n1441;
   wire n1442;
   wire n1443;
   wire n1444;
   wire n1445;
   wire n1446;
   wire n1447;
   wire n1448;
   wire n1449;
   wire n1450;
   wire n1451;
   wire n1452;
   wire n1453;
   wire n1454;
   wire n1455;
   wire n1456;
   wire n1457;
   wire n1458;
   wire n1459;
   wire n1460;
   wire n1461;
   wire n1462;
   wire n1463;
   wire n1464;
   wire n1465;
   wire n1466;
   wire n1467;
   wire n1468;
   wire n1469;
   wire n1470;
   wire n1471;
   wire n1472;
   wire n1473;
   wire n1474;
   wire n1475;
   wire n1476;
   wire n1477;
   wire n1478;
   wire n1479;
   wire n1480;
   wire n1481;
   wire n1482;
   wire n1483;
   wire n1484;
   wire n1485;
   wire n1486;
   wire n1487;
   wire n1488;
   wire n1489;
   wire n1490;
   wire n1491;
   wire n1492;
   wire n1493;
   wire n1494;
   wire n1495;
   wire n1496;
   wire n1497;
   wire n1498;
   wire n1499;
   wire n1500;
   wire n1501;
   wire n1502;
   wire n1503;
   wire n1504;
   wire n1505;
   wire n1506;
   wire n1507;
   wire n1508;
   wire n1509;
   wire n1510;
   wire n1511;
   wire n1512;
   wire n1513;
   wire n1514;
   wire n1515;
   wire n1516;
   wire n1517;
   wire n1518;
   wire n1519;
   wire n1520;
   wire n1521;
   wire n1522;
   wire n1523;
   wire n1524;
   wire n1525;
   wire n1526;
   wire n1527;
   wire n1528;
   wire n1529;
   wire n1530;
   wire n1531;
   wire n1532;
   wire n1533;
   wire n1534;
   wire n1535;
   wire n1536;
   wire n1537;
   wire n1538;
   wire n1539;
   wire n1540;
   wire n1541;
   wire n1542;
   wire n1543;
   wire n1544;
   wire n1545;
   wire n1546;
   wire n1547;
   wire n1548;
   wire n1549;
   wire n1550;
   wire n1551;
   wire n1552;
   wire n1553;
   wire n1554;
   wire n1555;
   wire n1556;
   wire n1557;
   wire n1558;
   wire n1559;
   wire n1560;
   wire n1561;
   wire n1562;
   wire n1563;
   wire n1564;
   wire n1565;
   wire n1566;
   wire n1567;
   wire n1568;
   wire n1569;
   wire n1570;
   wire n1571;
   wire n1572;
   wire n1573;
   wire n1574;
   wire n1575;
   wire n1576;
   wire n1577;
   wire n1578;
   wire n1579;
   wire n1580;
   wire n1581;
   wire n1582;
   wire n1583;
   wire n1584;
   wire n1585;
   wire n1586;
   wire n1587;
   wire n1588;
   wire n1589;
   wire n1590;
   wire n1591;
   wire n1592;
   wire n1593;
   wire n1594;
   wire n1595;
   wire n1596;
   wire n1597;
   wire n1598;
   wire n1599;
   wire n1600;
   wire n1601;
   wire n1602;
   wire n1603;
   wire n1604;
   wire n1605;
   wire n1606;
   wire n1607;
   wire n1608;
   wire n1609;
   wire n1610;
   wire n1611;
   wire n1612;
   wire n1613;
   wire n1614;
   wire n1615;
   wire n1616;
   wire n1617;
   wire n1618;
   wire n1619;
   wire n1620;
   wire n1621;
   wire n1622;
   wire n1623;
   wire n1624;
   wire n1625;
   wire n1626;
   wire n1627;
   wire n1628;
   wire n1629;
   wire n1630;
   wire n1631;
   wire n1632;
   wire n1633;
   wire n1634;
   wire n1635;
   wire n1636;
   wire n1637;
   wire n1638;
   wire n1639;
   wire n1640;
   wire n1641;
   wire n1642;
   wire n1643;
   wire n1644;
   wire n1645;
   wire n1646;
   wire n1647;
   wire n1648;
   wire n1649;
   wire n1650;
   wire n1651;
   wire n1652;
   wire n1653;
   wire n1654;
   wire n1655;
   wire n1656;
   wire n1657;
   wire n1658;
   wire n1659;
   wire n1660;
   wire n1661;
   wire n1662;
   wire n1663;
   wire n1664;
   wire n1665;
   wire n1666;
   wire n1667;
   wire n1668;
   wire n1669;
   wire n1670;
   wire n1671;
   wire n1672;
   wire n1673;
   wire n1674;
   wire n1675;
   wire n1676;
   wire n1677;
   wire n1678;
   wire n1679;
   wire n1680;
   wire n1681;
   wire n1682;
   wire n1683;
   wire n1684;
   wire n1685;
   wire n1686;
   wire n1687;
   wire n1688;
   wire n1689;
   wire n1690;
   wire n1691;
   wire n1692;
   wire n1693;
   wire n1694;
   wire n1695;
   wire n1696;
   wire n1697;
   wire n1698;
   wire n1699;
   wire n1700;
   wire n1701;
   wire n1702;
   wire n1703;
   wire n1704;
   wire n1705;
   wire n1706;
   wire n1707;
   wire n1708;
   wire n1709;
   wire n1710;
   wire n1711;
   wire n1712;
   wire n1713;
   wire n1714;
   wire n1715;
   wire n1716;
   wire n1717;
   wire n1718;
   wire n1719;
   wire n1720;
   wire n1721;
   wire n1722;
   wire n1723;
   wire n1724;
   wire n1725;
   wire n1726;
   wire n1727;
   wire n1728;
   wire n1729;
   wire n1730;
   wire n1731;
   wire n1732;
   wire n1733;
   wire n1734;
   wire n1735;
   wire n1736;
   wire n1737;
   wire n1738;
   wire n1739;
   wire n1740;
   wire n1741;
   wire n1742;
   wire n1743;
   wire n1744;
   wire n1745;
   wire n1746;
   wire n1747;
   wire n1748;
   wire n1749;
   wire n1750;
   wire n1751;
   wire n1752;
   wire n1753;
   wire n1754;
   wire n1755;
   wire n1756;
   wire n1757;
   wire n1758;
   wire n1759;
   wire n1760;
   wire n1761;
   wire n1762;
   wire n1763;
   wire n1764;
   wire n1765;
   wire n1766;
   wire n1767;
   wire n1768;
   wire n1769;
   wire n1770;
   wire n1771;
   wire n1772;
   wire n1773;
   wire n1774;
   wire n1775;
   wire n1776;
   wire n1777;
   wire n1778;
   wire n1779;
   wire n1780;
   wire n1781;
   wire n1782;
   wire n1783;
   wire n1784;
   wire n1785;
   wire n1786;
   wire n1787;
   wire n1788;
   wire n1789;
   wire n1790;
   wire n1791;
   wire n1792;
   wire n1793;
   wire n1794;
   wire n1795;
   wire n1796;
   wire n1797;
   wire n1798;
   wire n1799;
   wire n1800;
   wire n1801;
   wire n1802;
   wire n1803;
   wire n1804;
   wire n1805;
   wire n1806;
   wire n1807;
   wire n1808;
   wire n1809;
   wire n1810;
   wire n1811;
   wire n1812;
   wire n1813;
   wire n1814;
   wire n1815;
   wire n1816;
   wire n1817;
   wire n1818;
   wire n1819;
   wire n1820;
   wire n1821;
   wire n1822;
   wire n1823;
   wire n1824;
   wire n1825;
   wire n1826;
   wire n1827;
   wire n1828;
   wire n1829;
   wire n1830;
   wire n1831;
   wire n1832;
   wire n1833;
   wire n1834;
   wire n1835;
   wire n1836;
   wire n1837;
   wire n1838;
   wire n1839;
   wire n1840;
   wire n1841;
   wire n1842;
   wire n1843;
   wire n1844;
   wire n1845;
   wire n1846;
   wire n1847;
   wire n1848;
   wire n1849;
   wire n1850;
   wire n1851;
   wire n1852;
   wire n1853;
   wire n1854;
   wire n1855;
   wire n1856;
   wire n1857;
   wire n1858;
   wire n1859;
   wire n1860;
   wire n1861;
   wire n1862;
   wire n1863;
   wire n1864;
   wire n1865;
   wire n1866;
   wire n1867;
   wire n1868;
   wire n1869;
   wire n1870;
   wire n1871;
   wire n1872;
   wire n1873;
   wire n1874;
   wire n1875;
   wire n1876;
   wire n1877;
   wire n1878;
   wire n1879;
   wire n1880;
   wire n1881;
   wire n1882;
   wire n1883;
   wire n1884;
   wire n1885;
   wire n1886;
   wire n1887;
   wire n1888;
   wire n1889;
   wire n1890;
   wire n1891;
   wire n1892;
   wire n1893;
   wire n1894;
   wire n1895;
   wire n1896;
   wire n1897;
   wire n1898;
   wire n1899;
   wire n1900;
   wire n1901;
   wire n1902;
   wire n1903;
   wire n1904;
   wire n1905;
   wire n1906;
   wire n1907;
   wire n1908;
   wire n1909;
   wire n1910;
   wire n1911;
   wire n1912;
   wire n1913;
   wire n1914;
   wire n1915;
   wire n1916;
   wire n1917;
   wire n1918;
   wire n1919;
   wire n1920;
   wire n1921;
   wire n1922;
   wire n1923;
   wire n1924;
   wire n1925;
   wire n1926;
   wire n1927;
   wire n1928;
   wire n1929;
   wire n1930;
   wire n1931;
   wire n1932;
   wire n1933;
   wire n1934;
   wire n1935;
   wire n1936;
   wire n1937;
   wire n1938;
   wire n1939;
   wire n1940;
   wire n1941;
   wire n1942;
   wire n1943;
   wire n1944;
   wire n1945;
   wire n1946;
   wire n1947;
   wire n1948;
   wire n1949;
   wire n1950;
   wire n1951;
   wire n1952;
   wire n1953;
   wire n1954;
   wire n1955;
   wire n1956;
   wire n1957;
   wire n1958;
   wire n1959;
   wire n1960;
   wire n1961;
   wire n1962;
   wire n1963;
   wire n1964;
   wire n1965;
   wire n1966;
   wire n1967;
   wire n1968;
   wire n1969;
   wire n1970;
   wire n1971;
   wire n1972;
   wire n1973;
   wire n1974;
   wire n1975;
   wire n1976;
   wire n1977;
   wire n1978;
   wire n1979;
   wire n1980;
   wire n1981;
   wire n1982;
   wire n1983;
   wire n1984;
   wire n1985;
   wire n1986;
   wire n1987;
   wire n1988;
   wire n1989;
   wire n1990;
   wire n1991;
   wire n1992;
   wire n1993;
   wire n1994;
   wire n1995;
   wire n1996;
   wire n1997;
   wire n1998;
   wire n1999;
   wire n2000;
   wire n2001;
   wire n2002;
   wire n2003;
   wire n2004;
   wire n2005;
   wire n2006;
   wire n2007;
   wire n2008;
   wire n2009;
   wire n2010;
   wire n2011;
   wire n2012;
   wire n2013;
   wire n2014;
   wire n2015;
   wire n2016;
   wire n2017;
   wire n2018;
   wire n2019;
   wire n2020;
   wire n2021;
   wire n2022;
   wire n2023;
   wire n2024;
   wire n2025;
   wire n2026;
   wire n2027;
   wire n2028;
   wire n2029;
   wire n2030;
   wire n2031;
   wire n2032;
   wire n2033;
   wire n2034;
   wire n2035;
   wire n2036;
   wire n2037;
   wire n2038;
   wire n2039;
   wire n2040;
   wire n2041;
   wire n2042;
   wire n2043;
   wire n2044;
   wire n2045;
   wire n2046;
   wire n2047;
   wire n2048;
   wire n2049;
   wire n2050;
   wire n2051;
   wire n2052;
   wire n2053;
   wire n2054;
   wire n2055;
   wire n2056;
   wire n2057;
   wire n2058;
   wire n2059;
   wire n2060;
   wire n2061;
   wire n2062;
   wire n2063;
   wire n2064;
   wire n2065;
   wire n2066;
   wire n2067;
   wire n2068;
   wire n2069;
   wire n2070;
   wire n2071;
   wire n2072;
   wire n2073;
   wire n2074;
   wire n2075;
   wire n2076;
   wire n2077;
   wire n2078;
   wire n2079;
   wire n2080;
   wire n2081;
   wire n2082;
   wire n2083;
   wire n2084;
   wire n2085;
   wire n2086;
   wire n2087;
   wire n2088;
   wire n2089;
   wire n2090;
   wire n2091;
   wire n2092;
   wire n2093;
   wire n2094;
   wire n2095;
   wire n2096;
   wire n2097;
   wire n2098;
   wire n2099;
   wire n2100;
   wire n2101;
   wire n2102;
   wire n2103;
   wire n2104;
   wire n2105;
   wire n2106;
   wire n2107;
   wire n2108;
   wire n2109;
   wire n2110;
   wire n2111;
   wire n2112;
   wire n2113;
   wire n2114;
   wire n2115;
   wire n2116;
   wire n2117;
   wire n2118;
   wire n2119;
   wire n2120;
   wire n2121;
   wire n2122;
   wire n2123;
   wire n2124;
   wire n2125;
   wire n2126;
   wire n2127;
   wire n2128;
   wire n2129;
   wire n2130;
   wire n1;
   wire n2;
   wire n3;
   wire n4;
   wire n5;
   wire n6;
   wire n7;
   wire n8;
   wire n9;
   wire n10;
   wire n11;
   wire n12;
   wire n13;
   wire n14;
   wire n15;
   wire n16;
   wire n17;
   wire n18;
   wire n19;
   wire n20;
   wire n21;
   wire n22;
   wire n23;
   wire n24;
   wire n25;
   wire n26;
   wire n27;
   wire n28;
   wire n29;
   wire n30;
   wire n31;
   wire n32;
   wire n33;
   wire n34;
   wire n35;
   wire n36;
   wire n37;
   wire n2131;
   wire n2132;
   wire n2133;
   wire n2134;
   wire n2135;
   wire n2136;
   wire n2137;
   wire n2138;
   wire n2139;
   wire n2140;
   wire n2141;
   wire n2142;
   wire n2143;
   wire n2144;
   wire n2145;
   wire n2146;
   wire n2147;
   wire n2148;
   wire n2149;
   wire n2150;
   wire n2151;
   wire n2152;
   wire n2153;
   wire n2154;
   wire n2155;
   wire n2156;
   wire n2157;
   wire n2158;
   wire n2159;
   wire n2160;
   wire n2161;
   wire n2162;
   wire n2163;
   wire n2164;
   wire n2165;
   wire n2166;
   wire n2167;
   wire n2168;
   wire n2169;
   wire n2170;
   wire n2171;
   wire n2172;
   wire n2173;
   wire n2174;
   wire n2175;
   wire n2176;
   wire n2177;
   wire n2178;
   wire n2179;
   wire n2180;
   wire n2181;
   wire n2182;
   wire n2183;
   wire n2184;
   wire n2185;
   wire n2186;
   wire n2187;
   wire n2188;
   wire n2189;
   wire n2190;
   wire n2191;
   wire n2192;
   wire n2193;
   wire n2194;
   wire n2195;
   wire n2196;
   wire n2197;
   wire n2198;
   wire n2199;
   wire n2200;
   wire n2201;
   wire n2202;
   wire n2203;
   wire n2204;
   wire n2205;
   wire n2206;
   wire n2207;
   wire n2208;
   wire n2209;
   wire n2210;
   wire n2211;
   wire n2212;
   wire n2213;
   wire n2214;
   wire n2215;
   wire n2216;
   wire n2217;
   wire n2218;
   wire n2219;
   wire n2220;
   wire n2221;
   wire n2222;
   wire n2223;
   wire n2224;
   wire n2225;
   wire n2226;
   wire n2227;
   wire n2228;
   wire n2229;
   wire n2230;
   wire n2231;
   wire n2232;
   wire n2233;
   wire n2234;
   wire n2235;
   wire n2236;
   wire n2237;
   wire n2238;
   wire n2239;
   wire n2240;
   wire n2241;
   wire n2242;
   wire n2243;
   wire n2244;
   wire n2245;
   wire n2246;
   wire n2247;
   wire n2248;
   wire n2249;
   wire n2250;
   wire n2251;
   wire n2252;
   wire n2253;
   wire n2254;
   wire n2255;
   wire n2256;
   wire n2257;
   wire n2258;
   wire n2259;
   wire n2260;
   wire n2261;
   wire n2262;
   wire n2263;
   wire n2264;
   wire n2265;
   wire n2266;
   wire n2267;
   wire n2268;
   wire n2269;
   wire n2270;
   wire n2271;
   wire n2272;
   wire n2273;
   wire n2274;
   wire n2275;
   wire n2276;
   wire n2277;
   wire n2278;
   wire n2279;
   wire n2280;
   wire n2281;
   wire n2282;
   wire n2283;
   wire n2284;
   wire n2285;
   wire n2286;
   wire n2287;
   wire n2288;
   wire n2289;
   wire n2290;
   wire n2291;
   wire n2292;
   wire n2293;
   wire n2294;
   wire n2295;
   wire n2296;
   wire n2297;
   wire n2298;
   wire n2299;
   wire n2300;
   wire n2301;
   wire n2302;
   wire n2303;
   wire n2304;
   wire n2305;
   wire n2306;
   wire n2307;
   wire n2308;
   wire n2309;
   wire n2310;
   wire n2311;
   wire n2312;
   wire n2313;
   wire n2314;
   wire n2315;
   wire n2316;
   wire n2317;
   wire n2318;
   wire n2319;
   wire n2320;
   wire n2321;
   wire n2322;
   wire n2323;
   wire n2324;
   wire n2325;
   wire n2326;
   wire n2327;
   wire n2328;
   wire n2329;
   wire n2330;
   wire n2331;
   wire n2332;
   wire n2333;
   wire n2334;
   wire n2335;
   wire n2336;
   wire n2337;
   wire n2338;
   wire n2339;
   wire n2340;
   wire n2341;
   wire n2342;
   wire n2343;
   wire n2344;
   wire n2345;
   wire n2346;
   wire n2347;
   wire n2348;
   wire n2349;
   wire n2350;
   wire n2351;
   wire n2352;
   wire n2353;
   wire n2354;
   wire n2355;
   wire n2356;
   wire n2357;
   wire n2358;
   wire n2359;
   wire n2360;
   wire n2361;
   wire n2362;
   wire n2363;
   wire n2364;
   wire n2365;
   wire n2366;
   wire n2367;
   wire n2368;
   wire n2369;
   wire n2370;
   wire n2371;
   wire n2372;
   wire n2373;
   wire n2374;
   wire n2375;
   wire n2376;
   wire n2377;
   wire n2378;
   wire n2379;
   wire n2380;
   wire n2381;
   wire n2382;
   wire n2383;
   wire n2384;
   wire n2385;
   wire n2386;
   wire n2387;
   wire n2388;
   wire n2389;
   wire n2390;
   wire n2391;
   wire n2392;
   wire n2393;
   wire n2394;
   wire n2395;
   wire n2396;
   wire n2397;
   wire n2398;
   wire n2399;
   wire n2400;
   wire n2401;
   wire n2402;
   wire n2403;
   wire n2404;
   wire n2405;
   wire n2406;
   wire n2407;
   wire n2408;
   wire n2409;
   wire n2410;
   wire n2411;
   wire n2412;
   wire n2413;
   wire n2414;
   wire n2415;
   wire n2416;
   wire n2417;
   wire n2418;
   wire n2419;
   wire n2420;
   wire n2421;
   wire n2422;
   wire n2423;
   wire n2424;
   wire n2425;
   wire n2426;
   wire n2427;
   wire n2428;
   wire n2429;
   wire n2430;
   wire n2431;
   wire n2432;
   wire n2433;
   wire n2434;
   wire n2435;
   wire n2436;
   wire n2437;
   wire n2438;
   wire n2439;
   wire n2440;
   wire n2441;
   wire n2442;
   wire n2443;
   wire n2444;
   wire n2445;
   wire n2446;
   wire n2447;
   wire n2448;
   wire n2449;
   wire n2450;
   wire n2451;
   wire n2452;
   wire n2453;
   wire n2454;
   wire n2455;
   wire n2456;
   wire n2457;
   wire n2458;
   wire n2459;
   wire n2460;
   wire n2461;
   wire n2462;
   wire n2463;
   wire n2464;
   wire n2465;
   wire n2466;
   wire n2467;
   wire n2468;
   wire n2469;
   wire n2470;
   wire n2471;
   wire n2472;
   wire n2473;
   wire n2474;
   wire n2475;
   wire n2476;
   wire n2477;
   wire n2478;
   wire n2479;
   wire n2480;
   wire n2481;
   wire n2482;
   wire n2483;
   wire n2484;
   wire n2485;
   wire n2486;
   wire n2487;
   wire n2488;
   wire n2489;
   wire n2490;
   wire n2491;
   wire n2492;
   wire n2493;
   wire n2494;
   wire n2495;
   wire n2496;
   wire n2497;
   wire n2498;
   wire n2499;
   wire n2500;
   wire n2501;
   wire n2502;
   wire n2503;
   wire n2504;
   wire n2505;
   wire n2506;
   wire n2507;
   wire n2508;
   wire n2509;
   wire n2510;
   wire n2511;
   wire n2512;
   wire n2513;
   wire n2514;
   wire n2515;
   wire n2516;
   wire n2517;
   wire n2518;
   wire n2519;
   wire n2520;
   wire n2521;
   wire n2522;
   wire n2523;
   wire n2524;
   wire n2525;
   wire n2526;
   wire n2527;
   wire n2528;
   wire n2529;
   wire n2530;
   wire n2531;
   wire n2532;
   wire n2533;
   wire n2534;
   wire n2535;
   wire n2536;
   wire n2537;
   wire n2538;
   wire n2539;
   wire n2540;
   wire n2541;
   wire n2542;
   wire n2543;
   wire n2544;
   wire n2545;
   wire n2546;
   wire n2547;
   wire n2548;
   wire n2549;
   wire n2550;
   wire n2551;
   wire n2552;
   wire n2553;
   wire n2554;
   wire n2555;
   wire n2556;
   wire n2557;
   wire n2558;
   wire n2559;
   wire n2560;
   wire n2561;
   wire n2562;
   wire n2563;
   wire n2564;
   wire n2565;
   wire n2566;
   wire n2567;
   wire n2568;
   wire n2569;
   wire n2570;
   wire n2571;
   wire n2572;
   wire n2573;
   wire n2574;
   wire n2575;
   wire n2576;
   wire n2577;
   wire n2578;
   wire n2579;
   wire n2580;
   wire n2581;
   wire n2582;
   wire n2583;
   wire n2584;
   wire n2585;
   wire n2586;
   wire n2587;
   wire n2588;
   wire n2589;
   wire n2590;
   wire n2591;
   wire n2592;
   wire n2593;
   wire n2594;
   wire n2595;
   wire n2596;
   wire n2597;
   wire n2598;
   wire n2599;
   wire n2600;
   wire n2601;
   wire n2602;
   wire n2603;
   wire n2604;
   wire n2605;
   wire n2606;
   wire n2607;
   wire n2608;
   wire n2609;
   wire n2610;
   wire n2611;
   wire n2612;
   wire n2613;
   wire n2614;
   wire n2615;
   wire n2616;
   wire n2617;
   wire n2618;
   wire n2619;
   wire n2620;
   wire n2621;
   wire n2622;
   wire n2623;
   wire n2624;
   wire n2625;
   wire n2626;
   wire n2627;
   wire n2628;
   wire n2629;
   wire n2630;
   wire n2631;
   wire n2632;
   wire n2633;
   wire n2634;
   wire n2635;
   wire n2636;
   wire n2637;
   wire n2638;
   wire n2639;
   wire n2640;
   wire n2641;
   wire n2642;
   wire n2643;
   wire n2644;
   wire n2645;
   wire n2646;
   wire n2647;
   wire n2648;
   wire n2649;
   wire n2650;
   wire n2651;
   wire n2652;
   wire n2653;
   wire n2654;
   wire n2655;
   wire n2656;
   wire n2657;
   wire n2658;
   wire n2659;
   wire n2660;
   wire n2661;
   wire n2662;
   wire n2663;
   wire n2664;
   wire n2665;
   wire n2666;
   wire n2667;
   wire n2668;
   wire n2669;
   wire n2670;
   wire n2671;
   wire n2672;
   wire n2673;
   wire n2674;
   wire n2675;
   wire n2676;
   wire n2677;
   wire n2678;
   wire n2679;
   wire n2680;
   wire n2681;
   wire n2682;
   wire n2683;
   wire n2684;
   wire n2685;
   wire n2686;
   wire n2687;
   wire n2688;
   wire n2689;
   wire n2690;
   wire n2691;
   wire n2692;
   wire n2693;
   wire n2694;
   wire n2695;
   wire n2696;
   wire n2697;
   wire n2698;
   wire n2699;
   wire n2700;
   wire n2701;
   wire n2702;
   wire n2703;
   wire n2704;
   wire n2705;
   wire n2706;
   wire n2707;
   wire n2708;
   wire n2709;
   wire n2710;
   wire n2711;
   wire n2712;
   wire n2713;
   wire n2714;
   wire n2715;
   wire n2716;
   wire n2717;
   wire n2718;
   wire n2719;
   wire n2720;
   wire n2721;
   wire n2722;
   wire n2723;
   wire n2724;
   wire n2725;
   wire n2726;
   wire n2727;
   wire n2728;
   wire n2729;
   wire n2730;
   wire n2731;
   wire n2732;
   wire n2733;
   wire n2734;
   wire n2735;
   wire n2736;
   wire n2737;
   wire n2738;
   wire n2739;
   wire n2740;
   wire n2741;
   wire n2742;
   wire n2743;
   wire n2744;
   wire n2745;
   wire n2746;
   wire n2747;
   wire n2748;
   wire n2749;
   wire n2750;
   wire n2751;
   wire n2752;
   wire n2753;
   wire n2754;
   wire n2755;
   wire n2756;
   wire n2757;
   wire n2758;
   wire n2759;
   wire n2760;
   wire n2761;
   wire n2762;
   wire n2763;
   wire n2764;
   wire n2765;
   wire n2766;
   wire n2767;
   wire n2768;
   wire n2769;
   wire n2770;
   wire n2771;
   wire n2772;
   wire n2773;
   wire n2774;
   wire n2775;
   wire n2776;
   wire n2777;
   wire n2778;
   wire n2779;
   wire n2780;
   wire n2781;
   wire n2782;
   wire n2783;
   wire n2784;
   wire n2785;
   wire n2902;
   wire n2903;
   wire n2904;
   wire n2905;
   wire n2906;
   wire n2907;
   wire n2908;
   wire n2909;
   wire n2910;
   wire n2911;
   wire n2912;
   wire n2913;
   wire n2914;
   wire n2915;
   wire n2916;
   wire n2917;
   wire n2918;
   wire n2919;
   wire n2920;
   wire n2921;
   wire n2922;
   wire n2923;
   wire n2924;
   wire n2925;
   wire n2926;
   wire n2927;
   wire n2928;
   wire n2929;
   wire n2930;
   wire n2931;
   wire n2932;
   wire n2933;
   wire n2934;
   wire n2935;
   wire n2936;
   wire n2937;
   wire n2938;
   wire n2939;
   wire n2940;
   wire n2941;
   wire n2942;
   wire n2943;
   wire n2944;
   wire n2945;
   wire n2946;
   wire n2947;
   wire n2948;
   wire n2949;
   wire n2950;
   wire n2951;
   wire n2952;
   wire n2953;
   wire n2954;
   wire n2955;
   wire n2956;
   wire n2957;
   wire n2958;
   wire n2959;
   wire n2960;
   wire n2961;
   wire n2962;
   wire n2963;
   wire n2964;
   wire n2965;
   wire n2966;
   wire n2967;
   wire n2968;
   wire n2969;
   wire n2970;
   wire n2971;
   wire n2972;
   wire n2973;
   wire n2974;
   wire n2975;
   wire n2976;
   wire n2977;
   wire n2978;
   wire n2979;
   wire n2980;
   wire n2981;
   wire n2982;
   wire n2983;
   wire n2984;
   wire n2985;
   wire n2986;
   wire n2987;
   wire n2988;
   wire n2989;
   wire n2990;
   wire n2991;
   wire n2992;
   wire n2993;
   wire n2994;
   wire n2995;
   wire n2996;
   wire n2997;
   wire n2998;
   wire n2999;
   wire n3000;
   wire n3001;
   wire n3002;
   wire n3003;
   wire n3004;
   wire n3005;
   wire n3006;
   wire n3007;
   wire n3008;
   wire n3009;
   wire n3010;
   wire n3011;
   wire n3012;
   wire n3013;
   wire n3014;
   wire n3015;
   wire n3016;
   wire n3017;
   wire n3018;
   wire n3019;
   wire n3020;
   wire n3021;
   wire n3022;
   wire n3023;
   wire n3024;
   wire n3025;
   wire n3026;
   wire n3027;
   wire n3028;
   wire n3029;
   wire n3030;
   wire n3031;
   wire n3032;
   wire n3033;
   wire n3034;
   wire n3035;
   wire n3036;
   wire n3037;
   wire n3038;
   wire n3039;
   wire n3040;
   wire n3041;
   wire n3042;
   wire n3043;
   wire n3044;
   wire n3045;
   wire n3046;
   wire n3047;
   wire n3048;
   wire n3049;
   wire n3050;
   wire n3051;
   wire n3052;
   wire n3053;
   wire n3054;
   wire n3055;
   wire n3056;
   wire n3057;
   wire n3058;
   wire n3059;
   wire n3060;
   wire n3061;
   wire n3062;
   wire n3063;
   wire n3064;
   wire n3065;
   wire n3066;
   wire n3067;
   wire n3068;
   wire n3069;
   wire n3070;
   wire n3071;
   wire n3072;
   wire n3073;
   wire n3074;
   wire n3075;
   wire n3076;
   wire n3077;
   wire n3078;
   wire n3079;
   wire n3080;
   wire n3081;
   wire n3082;
   wire n3083;
   wire n3084;
   wire n3085;
   wire n3086;
   wire n3087;
   wire n3088;
   wire n3089;
   wire n3090;
   wire n3091;
   wire n3092;
   wire n3093;
   wire n3094;
   wire n3095;
   wire n3096;
   wire n3097;
   wire n3098;
   wire n3099;
   wire n3100;
   wire n3101;
   wire n3102;
   wire n3103;
   wire n3104;
   wire n3105;
   wire n3106;
   wire n3107;
   wire n3108;
   wire n3109;
   wire n3110;
   wire n3111;
   wire n3112;
   wire n3113;
   wire n3114;
   wire n3115;
   wire n3116;
   wire n3117;
   wire n3118;
   wire n3119;
   wire n3120;
   wire n3121;
   wire n3122;
   wire n3123;
   wire n3124;
   wire n3125;
   wire n3126;
   wire n3127;
   wire n3128;
   wire n3129;
   wire n3130;
   wire n3131;
   wire n3132;
   wire n3133;
   wire n3134;
   wire n3135;
   wire n3136;
   wire n3137;
   wire n3138;
   wire n3139;
   wire n3140;
   wire n3141;
   wire n3142;
   wire n3143;
   wire n3144;
   wire n3145;
   wire n3146;
   wire n3147;
   wire n3148;
   wire n3149;
   wire n3150;
   wire n3151;
   wire n3152;
   wire n3153;
   wire n3154;
   wire n3155;
   wire n3156;
   wire n3157;
   wire n3158;
   wire n3159;
   wire n3160;
   wire n3161;
   wire n3162;
   wire n3163;
   wire n3164;
   wire n3165;
   wire n3166;
   wire n3167;
   wire n3168;
   wire n3169;
   wire n3170;
   wire n3171;
   wire n3172;
   wire n3173;
   wire n3174;
   wire n3175;
   wire n3176;
   wire n3177;
   wire n3178;
   wire n3179;
   wire n3180;
   wire n3181;
   wire n3182;
   wire n3183;
   wire n3184;
   wire n3185;
   wire n3186;
   wire n3187;
   wire n3188;
   wire n3189;
   wire n3190;
   wire n3191;
   wire n3192;
   wire n3193;
   wire n3194;
   wire n3195;
   wire n3196;
   wire n3197;
   wire n3198;
   wire n3199;
   wire n3200;
   wire n3201;
   wire n3202;
   wire n3203;
   wire n3204;
   wire n3205;
   wire n3206;
   wire n3207;
   wire n3208;
   wire n3209;
   wire n3210;
   wire n3211;
   wire n3212;
   wire n3213;
   wire n3214;
   wire n3215;
   wire n3216;
   wire n3217;
   wire n3218;
   wire n3219;
   wire n3220;
   wire n3221;
   wire n3222;
   wire n3223;
   wire n3224;
   wire n3225;
   wire n3226;
   wire n3227;
   wire n3228;
   wire n3229;
   wire n3230;
   wire n3231;
   wire n3232;
   wire n3233;
   wire n3234;
   wire n3235;
   wire n3236;
   wire n3237;
   wire n3238;
   wire n3239;
   wire n3240;
   wire n3241;
   wire n3242;
   wire n3243;
   wire n3244;
   wire n3245;
   wire n3246;
   wire n3247;
   wire n3248;
   wire n3249;
   wire n3250;
   wire n3251;
   wire n3252;
   wire n3253;
   wire n3254;
   wire n3255;
   wire n3256;
   wire n3257;
   wire n3258;
   wire n3259;
   wire n3260;
   wire n3261;
   wire n3262;
   wire n3263;
   wire n3264;
   wire n3265;
   wire n3266;
   wire n3267;
   wire n3268;
   wire n3269;
   wire n3270;
   wire n3271;
   wire n3272;
   wire n3273;
   wire n3274;
   wire n3275;
   wire n3276;
   wire n3277;
   wire n3278;
   wire n3279;
   wire n3280;
   wire n3281;
   wire n3282;
   wire n3283;
   wire n3284;
   wire n3285;
   wire n3286;
   wire n3287;
   wire n3288;
   wire n3289;
   wire n3290;
   wire n3291;
   wire n3292;
   wire n3293;
   wire n3294;
   wire n3295;
   wire n3296;
   wire n3297;
   wire n3298;
   wire n3299;
   wire n3300;
   wire n3301;
   wire n3302;
   wire n3303;
   wire n3304;
   wire n3305;
   wire n3306;
   wire n3307;
   wire n3308;
   wire n3309;
   wire n3310;
   wire n3311;
   wire n3312;
   wire n3313;
   wire n3314;
   wire n3315;
   wire n3316;
   wire n3317;
   wire n3318;
   wire n3319;
   wire n3320;
   wire n3321;
   wire n3322;
   wire n3323;
   wire n3324;
   wire n3325;
   wire n3326;
   wire n3327;
   wire n3328;
   wire n3329;
   wire n3330;
   wire n3331;
   wire n3332;
   wire n3333;
   wire n3334;
   wire n3335;
   wire n3336;
   wire n3337;
   wire n3338;
   wire n3339;
   wire n3340;
   wire n3341;
   wire n3342;
   wire n3343;
   wire n3344;
   wire n3345;
   wire n3346;
   wire n3347;
   wire n3348;
   wire n3349;
   wire n3350;
   wire n3351;
   wire n3352;
   wire n3353;
   wire n3354;
   wire n3355;
   wire n3356;
   wire n3357;
   wire n3358;
   wire n3359;
   wire n3360;
   wire n3361;
   wire n3362;
   wire n3363;
   wire n3364;
   wire n3365;
   wire n3366;
   wire n3367;
   wire n3368;
   wire n3369;
   wire n3370;
   wire n3371;
   wire n3372;
   wire n3373;
   wire n3374;
   wire n3375;
   wire n3376;
   wire n3377;
   wire n3378;
   wire n3379;
   wire n3380;
   wire n3381;
   wire n3382;
   wire n3383;
   wire n3384;
   wire n3385;
   wire n3386;
   wire n3387;
   wire n3388;
   wire n3389;
   wire n3390;
   wire n3391;
   wire n3392;
   wire n3393;
   wire n3394;
   wire n3395;
   wire n3396;
   wire n3397;
   wire n3398;
   wire n3399;
   wire n3400;
   wire n3401;
   wire n3402;
   wire n3403;
   wire n3404;
   wire n3405;
   wire n3406;
   wire n3407;
   wire n3408;
   wire n3409;
   wire n3410;
   wire n3411;
   wire n3412;
   wire n3413;
   wire n3414;
   wire n3415;
   wire n3416;
   wire n3417;
   wire n3418;
   wire n3419;
   wire n3420;
   wire n3421;
   wire n3422;
   wire n3423;
   wire n3424;
   wire n3425;
   wire n3426;
   wire n3427;
   wire n3428;
   wire n3429;
   wire n3430;
   wire n3431;
   wire n3432;
   wire n3433;
   wire n3434;
   wire n3435;
   wire n3436;
   wire n3437;
   wire n3438;
   wire n3439;
   wire n3440;
   wire n3441;
   wire n3442;
   wire n3443;
   wire n3444;
   wire n3445;
   wire n3446;
   wire n3447;
   wire n3448;
   wire n3449;
   wire n3450;
   wire n3451;
   wire n3452;
   wire n3453;
   wire n3454;
   wire n3455;
   wire n3456;
   wire n3457;
   wire n3458;
   wire n3459;
   wire n3460;
   wire n3461;
   wire n3462;
   wire n3463;
   wire n3464;
   wire n3465;
   wire n3466;
   wire n3467;
   wire n3468;
   wire n3469;
   wire n3470;
   wire n3471;
   wire n3472;
   wire n3473;
   wire n3474;
   wire n3475;
   wire n3476;
   wire n3477;
   wire n3478;
   wire n3479;
   wire n3480;
   wire n3481;
   wire n3482;
   wire n3483;
   wire n3484;
   wire n3485;
   wire n3486;
   wire n3487;
   wire n3488;
   wire n3489;
   wire n3490;
   wire n3491;
   wire n3492;
   wire n3493;
   wire n3494;
   wire n3495;
   wire n3496;
   wire n3497;
   wire n3498;
   wire n3499;
   wire n3500;
   wire n3501;
   wire n3502;
   wire n3503;
   wire n3504;
   wire n3505;
   wire n3506;
   wire n3507;
   wire n3508;
   wire n3509;
   wire n3510;
   wire n3511;
   wire n3512;
   wire n3513;
   wire n3514;
   wire n3515;
   wire n3516;
   wire n3517;
   wire n3518;
   wire n3519;
   wire n3520;
   wire n3521;
   wire n3522;
   wire n3523;
   wire n3524;
   wire n3525;
   wire n3526;
   wire n3527;
   wire n3528;
   wire n3529;
   wire n3530;
   wire n3531;
   wire n3532;
   wire n3533;
   wire n3534;
   wire n3535;
   wire n3536;
   wire n3537;
   wire n3538;
   wire n3539;
   wire n3540;
   wire n3541;
   wire n3542;
   wire n3543;
   wire n3544;
   wire n3545;
   wire n3546;
   wire n3547;
   wire n3548;
   wire n3549;
   wire n3550;
   wire n3551;
   wire n3552;
   wire n3553;
   wire n3554;
   wire n3555;
   wire n3556;
   wire n3557;
   wire n3558;
   wire n3559;
   wire n3560;
   wire n3561;
   wire n3562;
   wire n3563;
   wire n3564;
   wire n3565;
   wire n3566;
   wire n3567;
   wire n3568;
   wire n3569;
   wire n3570;
   wire n3571;
   wire n3572;
   wire n3573;
   wire n3574;
   wire n3575;
   wire n3576;
   wire n3577;
   wire n3578;
   wire n3579;
   wire n3580;
   wire n3581;
   wire n3582;
   wire n3583;
   wire n3584;
   wire n3585;
   wire n3586;
   wire n3587;
   wire n3588;
   wire n3589;
   wire n3590;
   wire n3591;
   wire n3592;
   wire n3593;
   wire n4005;
   wire n4006;
   wire n4007;
   wire n4008;
   wire n4009;
   wire n4010;
   wire n4011;
   wire n4012;
   wire n4013;
   wire n4014;
   wire n4015;
   wire n4016;
   wire n4017;
   wire n4018;
   wire n4019;
   wire n4020;
   wire n4021;
   wire n4022;
   wire n4023;
   wire n4024;
   wire n4025;
   wire n4026;
   wire n4027;
   wire n4028;
   wire n4029;
   wire n4030;
   wire n4031;
   wire n4032;
   wire n4033;
   wire n4034;
   wire n4035;
   wire n4036;
   wire n4037;
   wire n4038;
   wire n4039;
   wire n4040;
   wire n4041;
   wire [1023:0] REGISTERS;

   BUF_X2 FE_OFC136_n2761 (.A(n2761),
	.Z(FE_OFN136_n2761));
   CLKBUF_X3 FE_OFC135_n2761 (.A(n2761),
	.Z(FE_OFN135_n2761));
   CLKBUF_X3 FE_OFC134_n3573 (.A(FE_OFN133_n3573),
	.Z(FE_OFN134_n3573));
   CLKBUF_X3 FE_OFC133_n3573 (.A(n3573),
	.Z(FE_OFN133_n3573));
   CLKBUF_X3 FE_OFC132_n3570 (.A(n3570),
	.Z(FE_OFN132_n3570));
   CLKBUF_X3 FE_OFC131_n3570 (.A(n3570),
	.Z(FE_OFN131_n3570));
   CLKBUF_X3 FE_OFC114_n2768 (.A(n2768),
	.Z(FE_OFN114_n2768));
   CLKBUF_X3 FE_OFC113_n2768 (.A(n2768),
	.Z(FE_OFN113_n2768));
   BUF_X2 FE_OFC112_n2763 (.A(FE_OFN110_n2763),
	.Z(FE_OFN112_n2763));
   BUF_X1 FE_OFC111_n2763 (.A(n2763),
	.Z(FE_OFN111_n2763));
   BUF_X2 FE_OFC110_n2763 (.A(n2763),
	.Z(FE_OFN110_n2763));
   CLKBUF_X3 FE_OFC109_n3569 (.A(n3569),
	.Z(FE_OFN109_n3569));
   CLKBUF_X3 FE_OFC108_n3569 (.A(n3569),
	.Z(FE_OFN108_n3569));
   BUF_X2 FE_OFC107_n3576 (.A(FE_OFN105_n3576),
	.Z(FE_OFN107_n3576));
   BUF_X1 FE_OFC106_n3576 (.A(FE_OFN105_n3576),
	.Z(FE_OFN106_n3576));
   BUF_X2 FE_OFC105_n3576 (.A(n3576),
	.Z(FE_OFN105_n3576));
   BUF_X2 FE_OFC89_n4027 (.A(n4027),
	.Z(FE_OFN89_n4027));
   BUF_X2 FE_OFC88_n4010 (.A(n4010),
	.Z(FE_OFN88_n4010));
   BUF_X2 FE_OFC87_n4032 (.A(n4032),
	.Z(FE_OFN87_n4032));
   BUF_X2 FE_OFC86_n4008 (.A(n4008),
	.Z(FE_OFN86_n4008));
   BUF_X2 FE_OFC85_n4022 (.A(n4022),
	.Z(FE_OFN85_n4022));
   BUF_X2 FE_OFC84_n4005 (.A(n4005),
	.Z(FE_OFN84_n4005));
   BUF_X2 FE_OFC83_n4024 (.A(n4024),
	.Z(FE_OFN83_n4024));
   BUF_X2 FE_OFC82_n4007 (.A(n4007),
	.Z(FE_OFN82_n4007));
   BUF_X2 FE_OFC81_n4030 (.A(n4030),
	.Z(FE_OFN81_n4030));
   BUF_X2 FE_OFC80_n4035 (.A(n4035),
	.Z(FE_OFN80_n4035));
   BUF_X2 FE_OFC79_n4023 (.A(n4023),
	.Z(FE_OFN79_n4023));
   BUF_X2 FE_OFC78_n4014 (.A(n4014),
	.Z(FE_OFN78_n4014));
   BUF_X2 FE_OFC77_n4026 (.A(n4026),
	.Z(FE_OFN77_n4026));
   BUF_X2 FE_OFC76_n4013 (.A(n4013),
	.Z(FE_OFN76_n4013));
   BUF_X2 FE_OFC75_n4028 (.A(n4028),
	.Z(FE_OFN75_n4028));
   BUF_X2 FE_OFC74_n4015 (.A(n4015),
	.Z(FE_OFN74_n4015));
   BUF_X2 FE_OFC73_n4009 (.A(n4009),
	.Z(FE_OFN73_n4009));
   BUF_X2 FE_OFC72_n4021 (.A(n4021),
	.Z(FE_OFN72_n4021));
   CLKBUF_X3 FE_OFC71_n4006 (.A(n4006),
	.Z(FE_OFN71_n4006));
   CLKBUF_X3 FE_OFC70_n4033 (.A(n4033),
	.Z(FE_OFN70_n4033));
   CLKBUF_X3 FE_OFC69_n4025 (.A(n4025),
	.Z(FE_OFN69_n4025));
   BUF_X2 FE_OFC68_n4011 (.A(n4011),
	.Z(FE_OFN68_n4011));
   BUF_X2 FE_OFC67_n4029 (.A(n4029),
	.Z(FE_OFN67_n4029));
   CLKBUF_X3 FE_OFC66_n4017 (.A(n4017),
	.Z(FE_OFN66_n4017));
   CLKBUF_X3 FE_OFC65_n4018 (.A(n4018),
	.Z(FE_OFN65_n4018));
   BUF_X2 FE_OFC64_n4012 (.A(n4012),
	.Z(FE_OFN64_n4012));
   CLKBUF_X3 FE_OFC63_n4031 (.A(n4031),
	.Z(FE_OFN63_n4031));
   CLKBUF_X3 FE_OFC62_n4016 (.A(n4016),
	.Z(FE_OFN62_n4016));
   BUF_X2 FE_OFC61_n4019 (.A(n4019),
	.Z(FE_OFN61_n4019));
   BUF_X2 FE_OFC60_n4036 (.A(n4036),
	.Z(FE_OFN60_n4036));
   CLKBUF_X3 FE_OFC59_n4034 (.A(n4034),
	.Z(FE_OFN59_n4034));
   BUF_X1 FE_OFC56_n2764 (.A(FE_OFN55_n2764),
	.Z(FE_OFN56_n2764));
   BUF_X2 FE_OFC55_n2764 (.A(FE_OFN54_n2764),
	.Z(FE_OFN55_n2764));
   CLKBUF_X3 FE_OFC54_n2764 (.A(n2764),
	.Z(FE_OFN54_n2764));
   BUF_X2 FE_OFC53_n2765 (.A(FE_OFN52_n2765),
	.Z(FE_OFN53_n2765));
   BUF_X1 FE_OFC52_n2765 (.A(n2765),
	.Z(FE_OFN52_n2765));
   BUF_X2 FE_OFC51_n2765 (.A(n2765),
	.Z(FE_OFN51_n2765));
   BUF_X1 FE_OFC50_n3575 (.A(FE_OFN49_n3575),
	.Z(FE_OFN50_n3575));
   BUF_X2 FE_OFC49_n3575 (.A(FE_OFN48_n3575),
	.Z(FE_OFN49_n3575));
   BUF_X2 FE_OFC48_n3575 (.A(n3575),
	.Z(FE_OFN48_n3575));
   CLKBUF_X3 FE_OFC47_n3572 (.A(FE_OFN46_n3572),
	.Z(FE_OFN47_n3572));
   CLKBUF_X3 FE_OFC46_n3572 (.A(n3572),
	.Z(FE_OFN46_n3572));
   BUF_X2 FE_OFC38_n3588 (.A(n3588),
	.Z(FE_OFN38_n3588));
   BUF_X2 FE_OFC33_n3584 (.A(n3584),
	.Z(FE_OFN33_n3584));
   BUF_X2 FE_OFC32_n2776 (.A(n2776),
	.Z(FE_OFN32_n2776));
   BUF_X2 FE_OFC31_n3582 (.A(n3582),
	.Z(FE_OFN31_n3582));
   BUF_X2 FE_OFC30_n2774 (.A(n2774),
	.Z(FE_OFN30_n2774));
   BUF_X2 FE_OFC18_n4041 (.A(n4041),
	.Z(FE_OFN18_n4041));
   CLKBUF_X3 FE_OFC14_n2762 (.A(n2762),
	.Z(FE_OFN14_n2762));
   CLKBUF_X3 FE_OFC13_n2762 (.A(n2762),
	.Z(FE_OFN13_n2762));
   CLKBUF_X3 FE_OFC12_n2767 (.A(FE_OFN11_n2767),
	.Z(FE_OFN12_n2767));
   CLKBUF_X3 FE_OFC11_n2767 (.A(n2767),
	.Z(FE_OFN11_n2767));
   BUF_X1 FE_OFC10_n2766 (.A(FE_OFN9_n2766),
	.Z(FE_OFN10_n2766));
   CLKBUF_X3 FE_OFC9_n2766 (.A(FE_OFN8_n2766),
	.Z(FE_OFN9_n2766));
   CLKBUF_X3 FE_OFC8_n2766 (.A(n2766),
	.Z(FE_OFN8_n2766));
   CLKBUF_X3 FE_OFC7_n3571 (.A(FE_OFN6_n3571),
	.Z(FE_OFN7_n3571));
   CLKBUF_X3 FE_OFC6_n3571 (.A(n3571),
	.Z(FE_OFN6_n3571));
   BUF_X2 FE_OFC5_n3574 (.A(FE_OFN4_n3574),
	.Z(FE_OFN5_n3574));
   BUF_X2 FE_OFC4_n3574 (.A(FE_OFN3_n3574),
	.Z(FE_OFN4_n3574));
   BUF_X1 FE_OFC3_n3574 (.A(n3574),
	.Z(FE_OFN3_n3574));
   DFF_X1 REGISTERS_reg_0__31_ (.D(n2130),
	.CK(CLK),
	.Q(REGISTERS[1023]));
   DFF_X1 REGISTERS_reg_0__30_ (.D(n2129),
	.CK(CLK),
	.Q(REGISTERS[1022]));
   DFF_X1 REGISTERS_reg_0__29_ (.D(n2128),
	.CK(CLK),
	.Q(REGISTERS[1021]));
   DFF_X1 REGISTERS_reg_0__28_ (.D(n2127),
	.CK(CLK),
	.Q(REGISTERS[1020]));
   DFF_X1 REGISTERS_reg_0__27_ (.D(n2126),
	.CK(CLK),
	.Q(REGISTERS[1019]));
   DFF_X1 REGISTERS_reg_0__26_ (.D(n2125),
	.CK(CLK),
	.Q(REGISTERS[1018]));
   DFF_X1 REGISTERS_reg_0__25_ (.D(n2124),
	.CK(CLK),
	.Q(REGISTERS[1017]));
   DFF_X1 REGISTERS_reg_0__24_ (.D(n2123),
	.CK(CLK),
	.Q(REGISTERS[1016]));
   DFF_X1 REGISTERS_reg_0__23_ (.D(n2122),
	.CK(CLK),
	.Q(REGISTERS[1015]));
   DFF_X1 REGISTERS_reg_0__22_ (.D(n2121),
	.CK(CLK),
	.Q(REGISTERS[1014]));
   DFF_X1 REGISTERS_reg_0__21_ (.D(n2120),
	.CK(CLK),
	.Q(REGISTERS[1013]));
   DFF_X1 REGISTERS_reg_0__20_ (.D(n2119),
	.CK(CLK),
	.Q(REGISTERS[1012]));
   DFF_X1 REGISTERS_reg_0__19_ (.D(n2118),
	.CK(CLK),
	.Q(REGISTERS[1011]));
   DFF_X1 REGISTERS_reg_0__18_ (.D(n2117),
	.CK(CLK),
	.Q(REGISTERS[1010]));
   DFF_X1 REGISTERS_reg_0__17_ (.D(n2116),
	.CK(CLK),
	.Q(REGISTERS[1009]));
   DFF_X1 REGISTERS_reg_0__16_ (.D(n2115),
	.CK(CLK),
	.Q(REGISTERS[1008]));
   DFF_X1 REGISTERS_reg_0__15_ (.D(n2114),
	.CK(CLK),
	.Q(REGISTERS[1007]));
   DFF_X1 REGISTERS_reg_0__14_ (.D(n2113),
	.CK(CLK),
	.Q(REGISTERS[1006]));
   DFF_X1 REGISTERS_reg_0__13_ (.D(n2112),
	.CK(CLK),
	.Q(REGISTERS[1005]));
   DFF_X1 REGISTERS_reg_0__12_ (.D(n2111),
	.CK(CLK),
	.Q(REGISTERS[1004]));
   DFF_X1 REGISTERS_reg_0__11_ (.D(n2110),
	.CK(CLK),
	.Q(REGISTERS[1003]));
   DFF_X1 REGISTERS_reg_0__10_ (.D(n2109),
	.CK(CLK),
	.Q(REGISTERS[1002]));
   DFF_X1 REGISTERS_reg_0__9_ (.D(n2108),
	.CK(CLK),
	.Q(REGISTERS[1001]));
   DFF_X1 REGISTERS_reg_0__8_ (.D(n2107),
	.CK(CLK),
	.Q(REGISTERS[1000]));
   DFF_X1 REGISTERS_reg_0__7_ (.D(n2106),
	.CK(CLK),
	.Q(REGISTERS[999]));
   DFF_X1 REGISTERS_reg_0__6_ (.D(n2105),
	.CK(CLK),
	.Q(REGISTERS[998]));
   DFF_X1 REGISTERS_reg_0__5_ (.D(n2104),
	.CK(CLK),
	.Q(REGISTERS[997]));
   DFF_X1 REGISTERS_reg_0__4_ (.D(n2103),
	.CK(CLK),
	.Q(REGISTERS[996]));
   DFF_X1 REGISTERS_reg_0__3_ (.D(n2102),
	.CK(CLK),
	.Q(REGISTERS[995]));
   DFF_X1 REGISTERS_reg_0__2_ (.D(n2101),
	.CK(CLK),
	.Q(REGISTERS[994]));
   DFF_X1 REGISTERS_reg_0__1_ (.D(n2100),
	.CK(CLK),
	.Q(REGISTERS[993]));
   DFF_X1 REGISTERS_reg_0__0_ (.D(n2099),
	.CK(CLK),
	.Q(REGISTERS[992]));
   DFF_X1 REGISTERS_reg_1__31_ (.D(n2098),
	.CK(CLK),
	.Q(REGISTERS[991]));
   DFF_X1 REGISTERS_reg_1__30_ (.D(n2097),
	.CK(CLK),
	.Q(REGISTERS[990]));
   DFF_X1 REGISTERS_reg_1__29_ (.D(n2096),
	.CK(CLK),
	.Q(REGISTERS[989]));
   DFF_X1 REGISTERS_reg_1__28_ (.D(n2095),
	.CK(CLK),
	.Q(REGISTERS[988]));
   DFF_X1 REGISTERS_reg_1__27_ (.D(n2094),
	.CK(CLK),
	.Q(REGISTERS[987]));
   DFF_X1 REGISTERS_reg_1__26_ (.D(n2093),
	.CK(CLK),
	.Q(REGISTERS[986]));
   DFF_X1 REGISTERS_reg_1__25_ (.D(n2092),
	.CK(CLK),
	.Q(REGISTERS[985]));
   DFF_X1 REGISTERS_reg_1__24_ (.D(n2091),
	.CK(CLK),
	.Q(REGISTERS[984]));
   DFF_X1 REGISTERS_reg_1__23_ (.D(n2090),
	.CK(CLK),
	.Q(REGISTERS[983]));
   DFF_X1 REGISTERS_reg_1__22_ (.D(n2089),
	.CK(CLK),
	.Q(REGISTERS[982]));
   DFF_X1 REGISTERS_reg_1__21_ (.D(n2088),
	.CK(CLK),
	.Q(REGISTERS[981]));
   DFF_X1 REGISTERS_reg_1__20_ (.D(n2087),
	.CK(CLK),
	.Q(REGISTERS[980]));
   DFF_X1 REGISTERS_reg_1__19_ (.D(n2086),
	.CK(CLK),
	.Q(REGISTERS[979]));
   DFF_X1 REGISTERS_reg_1__18_ (.D(n2085),
	.CK(CLK),
	.Q(REGISTERS[978]));
   DFF_X1 REGISTERS_reg_1__17_ (.D(n2084),
	.CK(CLK),
	.Q(REGISTERS[977]));
   DFF_X1 REGISTERS_reg_1__16_ (.D(n2083),
	.CK(CLK),
	.Q(REGISTERS[976]));
   DFF_X1 REGISTERS_reg_1__15_ (.D(n2082),
	.CK(CLK),
	.Q(REGISTERS[975]));
   DFF_X1 REGISTERS_reg_1__14_ (.D(n2081),
	.CK(CLK),
	.Q(REGISTERS[974]));
   DFF_X1 REGISTERS_reg_1__13_ (.D(n2080),
	.CK(CLK),
	.Q(REGISTERS[973]));
   DFF_X1 REGISTERS_reg_1__12_ (.D(n2079),
	.CK(CLK),
	.Q(REGISTERS[972]));
   DFF_X1 REGISTERS_reg_1__11_ (.D(n2078),
	.CK(CLK),
	.Q(REGISTERS[971]));
   DFF_X1 REGISTERS_reg_1__10_ (.D(n2077),
	.CK(CLK),
	.Q(REGISTERS[970]));
   DFF_X1 REGISTERS_reg_1__9_ (.D(n2076),
	.CK(CLK),
	.Q(REGISTERS[969]));
   DFF_X1 REGISTERS_reg_1__8_ (.D(n2075),
	.CK(CLK),
	.Q(REGISTERS[968]));
   DFF_X1 REGISTERS_reg_1__7_ (.D(n2074),
	.CK(CLK),
	.Q(REGISTERS[967]));
   DFF_X1 REGISTERS_reg_1__6_ (.D(n2073),
	.CK(CLK),
	.Q(REGISTERS[966]));
   DFF_X1 REGISTERS_reg_1__5_ (.D(n2072),
	.CK(CLK),
	.Q(REGISTERS[965]));
   DFF_X1 REGISTERS_reg_1__4_ (.D(n2071),
	.CK(CLK),
	.Q(REGISTERS[964]));
   DFF_X1 REGISTERS_reg_1__3_ (.D(n2070),
	.CK(CLK),
	.Q(REGISTERS[963]));
   DFF_X1 REGISTERS_reg_1__2_ (.D(n2069),
	.CK(CLK),
	.Q(REGISTERS[962]));
   DFF_X1 REGISTERS_reg_1__1_ (.D(n2068),
	.CK(CLK),
	.Q(REGISTERS[961]));
   DFF_X1 REGISTERS_reg_1__0_ (.D(n2067),
	.CK(CLK),
	.Q(REGISTERS[960]));
   DFF_X1 REGISTERS_reg_2__31_ (.D(n2066),
	.CK(CLK),
	.Q(REGISTERS[959]));
   DFF_X1 REGISTERS_reg_2__30_ (.D(n2065),
	.CK(CLK),
	.Q(REGISTERS[958]));
   DFF_X1 REGISTERS_reg_2__29_ (.D(n2064),
	.CK(CLK),
	.Q(REGISTERS[957]));
   DFF_X1 REGISTERS_reg_2__28_ (.D(n2063),
	.CK(CLK),
	.Q(REGISTERS[956]));
   DFF_X1 REGISTERS_reg_2__27_ (.D(n2062),
	.CK(CLK),
	.Q(REGISTERS[955]));
   DFF_X1 REGISTERS_reg_2__26_ (.D(n2061),
	.CK(CLK),
	.Q(REGISTERS[954]));
   DFF_X1 REGISTERS_reg_2__25_ (.D(n2060),
	.CK(CLK),
	.Q(REGISTERS[953]));
   DFF_X1 REGISTERS_reg_2__24_ (.D(n2059),
	.CK(CLK),
	.Q(REGISTERS[952]));
   DFF_X1 REGISTERS_reg_2__23_ (.D(n2058),
	.CK(CLK),
	.Q(REGISTERS[951]));
   DFF_X1 REGISTERS_reg_2__22_ (.D(n2057),
	.CK(CLK),
	.Q(REGISTERS[950]));
   DFF_X1 REGISTERS_reg_2__21_ (.D(n2056),
	.CK(CLK),
	.Q(REGISTERS[949]));
   DFF_X1 REGISTERS_reg_2__20_ (.D(n2055),
	.CK(CLK),
	.Q(REGISTERS[948]));
   DFF_X1 REGISTERS_reg_2__19_ (.D(n2054),
	.CK(CLK),
	.Q(REGISTERS[947]));
   DFF_X1 REGISTERS_reg_2__18_ (.D(n2053),
	.CK(CLK),
	.Q(REGISTERS[946]));
   DFF_X1 REGISTERS_reg_2__17_ (.D(n2052),
	.CK(CLK),
	.Q(REGISTERS[945]));
   DFF_X1 REGISTERS_reg_2__16_ (.D(n2051),
	.CK(CLK),
	.Q(REGISTERS[944]));
   DFF_X1 REGISTERS_reg_2__15_ (.D(n2050),
	.CK(CLK),
	.Q(REGISTERS[943]));
   DFF_X1 REGISTERS_reg_2__14_ (.D(n2049),
	.CK(CLK),
	.Q(REGISTERS[942]));
   DFF_X1 REGISTERS_reg_2__13_ (.D(n2048),
	.CK(CLK),
	.Q(REGISTERS[941]));
   DFF_X1 REGISTERS_reg_2__12_ (.D(n2047),
	.CK(CLK),
	.Q(REGISTERS[940]));
   DFF_X1 REGISTERS_reg_2__11_ (.D(n2046),
	.CK(CLK),
	.Q(REGISTERS[939]));
   DFF_X1 REGISTERS_reg_2__10_ (.D(n2045),
	.CK(CLK),
	.Q(REGISTERS[938]));
   DFF_X1 REGISTERS_reg_2__9_ (.D(n2044),
	.CK(CLK),
	.Q(REGISTERS[937]));
   DFF_X1 REGISTERS_reg_2__8_ (.D(n2043),
	.CK(CLK),
	.Q(REGISTERS[936]));
   DFF_X1 REGISTERS_reg_2__7_ (.D(n2042),
	.CK(CLK),
	.Q(REGISTERS[935]));
   DFF_X1 REGISTERS_reg_2__6_ (.D(n2041),
	.CK(CLK),
	.Q(REGISTERS[934]));
   DFF_X1 REGISTERS_reg_2__5_ (.D(n2040),
	.CK(CLK),
	.Q(REGISTERS[933]));
   DFF_X1 REGISTERS_reg_2__4_ (.D(n2039),
	.CK(CLK),
	.Q(REGISTERS[932]));
   DFF_X1 REGISTERS_reg_2__3_ (.D(n2038),
	.CK(CLK),
	.Q(REGISTERS[931]));
   DFF_X1 REGISTERS_reg_2__2_ (.D(n2037),
	.CK(CLK),
	.Q(REGISTERS[930]));
   DFF_X1 REGISTERS_reg_2__1_ (.D(n2036),
	.CK(CLK),
	.Q(REGISTERS[929]));
   DFF_X1 REGISTERS_reg_2__0_ (.D(n2035),
	.CK(CLK),
	.Q(REGISTERS[928]));
   DFF_X1 REGISTERS_reg_3__31_ (.D(n2034),
	.CK(CLK),
	.Q(REGISTERS[927]));
   DFF_X1 REGISTERS_reg_3__30_ (.D(n2033),
	.CK(CLK),
	.Q(REGISTERS[926]));
   DFF_X1 REGISTERS_reg_3__29_ (.D(n2032),
	.CK(CLK),
	.Q(REGISTERS[925]));
   DFF_X1 REGISTERS_reg_3__28_ (.D(n2031),
	.CK(CLK),
	.Q(REGISTERS[924]));
   DFF_X1 REGISTERS_reg_3__27_ (.D(n2030),
	.CK(CLK),
	.Q(REGISTERS[923]));
   DFF_X1 REGISTERS_reg_3__26_ (.D(n2029),
	.CK(CLK),
	.Q(REGISTERS[922]));
   DFF_X1 REGISTERS_reg_3__25_ (.D(n2028),
	.CK(CLK),
	.Q(REGISTERS[921]));
   DFF_X1 REGISTERS_reg_3__24_ (.D(n2027),
	.CK(CLK),
	.Q(REGISTERS[920]));
   DFF_X1 REGISTERS_reg_3__23_ (.D(n2026),
	.CK(CLK),
	.Q(REGISTERS[919]));
   DFF_X1 REGISTERS_reg_3__22_ (.D(n2025),
	.CK(CLK),
	.Q(REGISTERS[918]));
   DFF_X1 REGISTERS_reg_3__21_ (.D(n2024),
	.CK(CLK),
	.Q(REGISTERS[917]));
   DFF_X1 REGISTERS_reg_3__20_ (.D(n2023),
	.CK(CLK),
	.Q(REGISTERS[916]));
   DFF_X1 REGISTERS_reg_3__19_ (.D(n2022),
	.CK(CLK),
	.Q(REGISTERS[915]));
   DFF_X1 REGISTERS_reg_3__18_ (.D(n2021),
	.CK(CLK),
	.Q(REGISTERS[914]));
   DFF_X1 REGISTERS_reg_3__17_ (.D(n2020),
	.CK(CLK),
	.Q(REGISTERS[913]));
   DFF_X1 REGISTERS_reg_3__16_ (.D(n2019),
	.CK(CLK),
	.Q(REGISTERS[912]));
   DFF_X1 REGISTERS_reg_3__15_ (.D(n2018),
	.CK(CLK),
	.Q(REGISTERS[911]));
   DFF_X1 REGISTERS_reg_3__14_ (.D(n2017),
	.CK(CLK),
	.Q(REGISTERS[910]));
   DFF_X1 REGISTERS_reg_3__13_ (.D(n2016),
	.CK(CLK),
	.Q(REGISTERS[909]));
   DFF_X1 REGISTERS_reg_3__12_ (.D(n2015),
	.CK(CLK),
	.Q(REGISTERS[908]));
   DFF_X1 REGISTERS_reg_3__11_ (.D(n2014),
	.CK(CLK),
	.Q(REGISTERS[907]));
   DFF_X1 REGISTERS_reg_3__10_ (.D(n2013),
	.CK(CLK),
	.Q(REGISTERS[906]));
   DFF_X1 REGISTERS_reg_3__9_ (.D(n2012),
	.CK(CLK),
	.Q(REGISTERS[905]));
   DFF_X1 REGISTERS_reg_3__8_ (.D(n2011),
	.CK(CLK),
	.Q(REGISTERS[904]));
   DFF_X1 REGISTERS_reg_3__7_ (.D(n2010),
	.CK(CLK),
	.Q(REGISTERS[903]));
   DFF_X1 REGISTERS_reg_3__6_ (.D(n2009),
	.CK(CLK),
	.Q(REGISTERS[902]));
   DFF_X1 REGISTERS_reg_3__5_ (.D(n2008),
	.CK(CLK),
	.Q(REGISTERS[901]));
   DFF_X1 REGISTERS_reg_3__4_ (.D(n2007),
	.CK(CLK),
	.Q(REGISTERS[900]));
   DFF_X1 REGISTERS_reg_3__3_ (.D(n2006),
	.CK(CLK),
	.Q(REGISTERS[899]));
   DFF_X1 REGISTERS_reg_3__2_ (.D(n2005),
	.CK(CLK),
	.Q(REGISTERS[898]));
   DFF_X1 REGISTERS_reg_3__1_ (.D(n2004),
	.CK(CLK),
	.Q(REGISTERS[897]));
   DFF_X1 REGISTERS_reg_3__0_ (.D(n2003),
	.CK(CLK),
	.Q(REGISTERS[896]));
   DFF_X1 REGISTERS_reg_4__31_ (.D(n2002),
	.CK(CLK),
	.Q(REGISTERS[895]));
   DFF_X1 REGISTERS_reg_4__30_ (.D(n2001),
	.CK(CLK),
	.Q(REGISTERS[894]));
   DFF_X1 REGISTERS_reg_4__29_ (.D(n2000),
	.CK(CLK),
	.Q(REGISTERS[893]));
   DFF_X1 REGISTERS_reg_4__28_ (.D(n1999),
	.CK(CLK),
	.Q(REGISTERS[892]));
   DFF_X1 REGISTERS_reg_4__27_ (.D(n1998),
	.CK(CLK),
	.Q(REGISTERS[891]));
   DFF_X1 REGISTERS_reg_4__26_ (.D(n1997),
	.CK(CLK),
	.Q(REGISTERS[890]));
   DFF_X1 REGISTERS_reg_4__25_ (.D(n1996),
	.CK(CLK),
	.Q(REGISTERS[889]));
   DFF_X1 REGISTERS_reg_4__24_ (.D(n1995),
	.CK(CLK),
	.Q(REGISTERS[888]));
   DFF_X1 REGISTERS_reg_4__23_ (.D(n1994),
	.CK(CLK),
	.Q(REGISTERS[887]));
   DFF_X1 REGISTERS_reg_4__22_ (.D(n1993),
	.CK(CLK),
	.Q(REGISTERS[886]));
   DFF_X1 REGISTERS_reg_4__21_ (.D(n1992),
	.CK(CLK),
	.Q(REGISTERS[885]));
   DFF_X1 REGISTERS_reg_4__20_ (.D(n1991),
	.CK(CLK),
	.Q(REGISTERS[884]));
   DFF_X1 REGISTERS_reg_4__19_ (.D(n1990),
	.CK(CLK),
	.Q(REGISTERS[883]));
   DFF_X1 REGISTERS_reg_4__18_ (.D(n1989),
	.CK(CLK),
	.Q(REGISTERS[882]));
   DFF_X1 REGISTERS_reg_4__17_ (.D(n1988),
	.CK(CLK),
	.Q(REGISTERS[881]));
   DFF_X1 REGISTERS_reg_4__16_ (.D(n1987),
	.CK(CLK),
	.Q(REGISTERS[880]));
   DFF_X1 REGISTERS_reg_4__15_ (.D(n1986),
	.CK(CLK),
	.Q(REGISTERS[879]));
   DFF_X1 REGISTERS_reg_4__14_ (.D(n1985),
	.CK(CLK),
	.Q(REGISTERS[878]));
   DFF_X1 REGISTERS_reg_4__13_ (.D(n1984),
	.CK(CLK),
	.Q(REGISTERS[877]));
   DFF_X1 REGISTERS_reg_4__12_ (.D(n1983),
	.CK(CLK),
	.Q(REGISTERS[876]));
   DFF_X1 REGISTERS_reg_4__11_ (.D(n1982),
	.CK(CLK),
	.Q(REGISTERS[875]));
   DFF_X1 REGISTERS_reg_4__10_ (.D(n1981),
	.CK(CLK),
	.Q(REGISTERS[874]));
   DFF_X1 REGISTERS_reg_4__9_ (.D(n1980),
	.CK(CLK),
	.Q(REGISTERS[873]));
   DFF_X1 REGISTERS_reg_4__8_ (.D(n1979),
	.CK(CLK),
	.Q(REGISTERS[872]));
   DFF_X1 REGISTERS_reg_4__7_ (.D(n1978),
	.CK(CLK),
	.Q(REGISTERS[871]));
   DFF_X1 REGISTERS_reg_4__6_ (.D(n1977),
	.CK(CLK),
	.Q(REGISTERS[870]));
   DFF_X1 REGISTERS_reg_4__5_ (.D(n1976),
	.CK(CLK),
	.Q(REGISTERS[869]));
   DFF_X1 REGISTERS_reg_4__4_ (.D(n1975),
	.CK(CLK),
	.Q(REGISTERS[868]));
   DFF_X1 REGISTERS_reg_4__3_ (.D(n1974),
	.CK(CLK),
	.Q(REGISTERS[867]));
   DFF_X1 REGISTERS_reg_4__2_ (.D(n1973),
	.CK(CLK),
	.Q(REGISTERS[866]));
   DFF_X1 REGISTERS_reg_4__1_ (.D(n1972),
	.CK(CLK),
	.Q(REGISTERS[865]));
   DFF_X1 REGISTERS_reg_4__0_ (.D(n1971),
	.CK(CLK),
	.Q(REGISTERS[864]));
   DFF_X1 REGISTERS_reg_5__31_ (.D(n1970),
	.CK(CLK),
	.Q(REGISTERS[863]));
   DFF_X1 REGISTERS_reg_5__30_ (.D(n1969),
	.CK(CLK),
	.Q(REGISTERS[862]));
   DFF_X1 REGISTERS_reg_5__29_ (.D(n1968),
	.CK(CLK),
	.Q(REGISTERS[861]));
   DFF_X1 REGISTERS_reg_5__28_ (.D(n1967),
	.CK(CLK),
	.Q(REGISTERS[860]));
   DFF_X1 REGISTERS_reg_5__27_ (.D(n1966),
	.CK(CLK),
	.Q(REGISTERS[859]));
   DFF_X1 REGISTERS_reg_5__26_ (.D(n1965),
	.CK(CLK),
	.Q(REGISTERS[858]));
   DFF_X1 REGISTERS_reg_5__25_ (.D(n1964),
	.CK(CLK),
	.Q(REGISTERS[857]));
   DFF_X1 REGISTERS_reg_5__24_ (.D(n1963),
	.CK(CLK),
	.Q(REGISTERS[856]));
   DFF_X1 REGISTERS_reg_5__23_ (.D(n1962),
	.CK(CLK),
	.Q(REGISTERS[855]));
   DFF_X1 REGISTERS_reg_5__22_ (.D(n1961),
	.CK(CLK),
	.Q(REGISTERS[854]));
   DFF_X1 REGISTERS_reg_5__21_ (.D(n1960),
	.CK(CLK),
	.Q(REGISTERS[853]));
   DFF_X1 REGISTERS_reg_5__20_ (.D(n1959),
	.CK(CLK),
	.Q(REGISTERS[852]));
   DFF_X1 REGISTERS_reg_5__19_ (.D(n1958),
	.CK(CLK),
	.Q(REGISTERS[851]));
   DFF_X1 REGISTERS_reg_5__18_ (.D(n1957),
	.CK(CLK),
	.Q(REGISTERS[850]));
   DFF_X1 REGISTERS_reg_5__17_ (.D(n1956),
	.CK(CLK),
	.Q(REGISTERS[849]));
   DFF_X1 REGISTERS_reg_5__16_ (.D(n1955),
	.CK(CLK),
	.Q(REGISTERS[848]));
   DFF_X1 REGISTERS_reg_5__15_ (.D(n1954),
	.CK(CLK),
	.Q(REGISTERS[847]));
   DFF_X1 REGISTERS_reg_5__14_ (.D(n1953),
	.CK(CLK),
	.Q(REGISTERS[846]));
   DFF_X1 REGISTERS_reg_5__13_ (.D(n1952),
	.CK(CLK),
	.Q(REGISTERS[845]));
   DFF_X1 REGISTERS_reg_5__12_ (.D(n1951),
	.CK(CLK),
	.Q(REGISTERS[844]));
   DFF_X1 REGISTERS_reg_5__11_ (.D(n1950),
	.CK(CLK),
	.Q(REGISTERS[843]));
   DFF_X1 REGISTERS_reg_5__10_ (.D(n1949),
	.CK(CLK),
	.Q(REGISTERS[842]));
   DFF_X1 REGISTERS_reg_5__9_ (.D(n1948),
	.CK(CLK),
	.Q(REGISTERS[841]));
   DFF_X1 REGISTERS_reg_5__8_ (.D(n1947),
	.CK(CLK),
	.Q(REGISTERS[840]));
   DFF_X1 REGISTERS_reg_5__7_ (.D(n1946),
	.CK(CLK),
	.Q(REGISTERS[839]));
   DFF_X1 REGISTERS_reg_5__6_ (.D(n1945),
	.CK(CLK),
	.Q(REGISTERS[838]));
   DFF_X1 REGISTERS_reg_5__5_ (.D(n1944),
	.CK(CLK),
	.Q(REGISTERS[837]));
   DFF_X1 REGISTERS_reg_5__4_ (.D(n1943),
	.CK(CLK),
	.Q(REGISTERS[836]));
   DFF_X1 REGISTERS_reg_5__3_ (.D(n1942),
	.CK(CLK),
	.Q(REGISTERS[835]));
   DFF_X1 REGISTERS_reg_5__2_ (.D(n1941),
	.CK(CLK),
	.Q(REGISTERS[834]));
   DFF_X1 REGISTERS_reg_5__1_ (.D(n1940),
	.CK(CLK),
	.Q(REGISTERS[833]));
   DFF_X1 REGISTERS_reg_5__0_ (.D(n1939),
	.CK(CLK),
	.Q(REGISTERS[832]));
   DFF_X1 REGISTERS_reg_6__31_ (.D(n1938),
	.CK(CLK),
	.Q(REGISTERS[831]));
   DFF_X1 REGISTERS_reg_6__30_ (.D(n1937),
	.CK(CLK),
	.Q(REGISTERS[830]));
   DFF_X1 REGISTERS_reg_6__29_ (.D(n1936),
	.CK(CLK),
	.Q(REGISTERS[829]));
   DFF_X1 REGISTERS_reg_6__28_ (.D(n1935),
	.CK(CLK),
	.Q(REGISTERS[828]));
   DFF_X1 REGISTERS_reg_6__27_ (.D(n1934),
	.CK(CLK),
	.Q(REGISTERS[827]));
   DFF_X1 REGISTERS_reg_6__26_ (.D(n1933),
	.CK(CLK),
	.Q(REGISTERS[826]));
   DFF_X1 REGISTERS_reg_6__25_ (.D(n1932),
	.CK(CLK),
	.Q(REGISTERS[825]));
   DFF_X1 REGISTERS_reg_6__24_ (.D(n1931),
	.CK(CLK),
	.Q(REGISTERS[824]));
   DFF_X1 REGISTERS_reg_6__23_ (.D(n1930),
	.CK(CLK),
	.Q(REGISTERS[823]));
   DFF_X1 REGISTERS_reg_6__22_ (.D(n1929),
	.CK(CLK),
	.Q(REGISTERS[822]));
   DFF_X1 REGISTERS_reg_6__21_ (.D(n1928),
	.CK(CLK),
	.Q(REGISTERS[821]));
   DFF_X1 REGISTERS_reg_6__20_ (.D(n1927),
	.CK(CLK),
	.Q(REGISTERS[820]));
   DFF_X1 REGISTERS_reg_6__19_ (.D(n1926),
	.CK(CLK),
	.Q(REGISTERS[819]));
   DFF_X1 REGISTERS_reg_6__18_ (.D(n1925),
	.CK(CLK),
	.Q(REGISTERS[818]));
   DFF_X1 REGISTERS_reg_6__17_ (.D(n1924),
	.CK(CLK),
	.Q(REGISTERS[817]));
   DFF_X1 REGISTERS_reg_6__16_ (.D(n1923),
	.CK(CLK),
	.Q(REGISTERS[816]));
   DFF_X1 REGISTERS_reg_6__15_ (.D(n1922),
	.CK(CLK),
	.Q(REGISTERS[815]));
   DFF_X1 REGISTERS_reg_6__14_ (.D(n1921),
	.CK(CLK),
	.Q(REGISTERS[814]));
   DFF_X1 REGISTERS_reg_6__13_ (.D(n1920),
	.CK(CLK),
	.Q(REGISTERS[813]));
   DFF_X1 REGISTERS_reg_6__12_ (.D(n1919),
	.CK(CLK),
	.Q(REGISTERS[812]));
   DFF_X1 REGISTERS_reg_6__11_ (.D(n1918),
	.CK(CLK),
	.Q(REGISTERS[811]));
   DFF_X1 REGISTERS_reg_6__10_ (.D(n1917),
	.CK(CLK),
	.Q(REGISTERS[810]));
   DFF_X1 REGISTERS_reg_6__9_ (.D(n1916),
	.CK(CLK),
	.Q(REGISTERS[809]));
   DFF_X1 REGISTERS_reg_6__8_ (.D(n1915),
	.CK(CLK),
	.Q(REGISTERS[808]));
   DFF_X1 REGISTERS_reg_6__7_ (.D(n1914),
	.CK(CLK),
	.Q(REGISTERS[807]));
   DFF_X1 REGISTERS_reg_6__6_ (.D(n1913),
	.CK(CLK),
	.Q(REGISTERS[806]));
   DFF_X1 REGISTERS_reg_6__5_ (.D(n1912),
	.CK(CLK),
	.Q(REGISTERS[805]));
   DFF_X1 REGISTERS_reg_6__4_ (.D(n1911),
	.CK(CLK),
	.Q(REGISTERS[804]));
   DFF_X1 REGISTERS_reg_6__3_ (.D(n1910),
	.CK(CLK),
	.Q(REGISTERS[803]));
   DFF_X1 REGISTERS_reg_6__2_ (.D(n1909),
	.CK(CLK),
	.Q(REGISTERS[802]));
   DFF_X1 REGISTERS_reg_6__1_ (.D(n1908),
	.CK(CLK),
	.Q(REGISTERS[801]));
   DFF_X1 REGISTERS_reg_6__0_ (.D(n1907),
	.CK(CLK),
	.Q(REGISTERS[800]));
   DFF_X1 REGISTERS_reg_7__31_ (.D(n1906),
	.CK(CLK),
	.Q(REGISTERS[799]));
   DFF_X1 REGISTERS_reg_7__30_ (.D(n1905),
	.CK(CLK),
	.Q(REGISTERS[798]));
   DFF_X1 REGISTERS_reg_7__29_ (.D(n1904),
	.CK(CLK),
	.Q(REGISTERS[797]));
   DFF_X1 REGISTERS_reg_7__28_ (.D(n1903),
	.CK(CLK),
	.Q(REGISTERS[796]));
   DFF_X1 REGISTERS_reg_7__27_ (.D(n1902),
	.CK(CLK),
	.Q(REGISTERS[795]));
   DFF_X1 REGISTERS_reg_7__26_ (.D(n1901),
	.CK(CLK),
	.Q(REGISTERS[794]));
   DFF_X1 REGISTERS_reg_7__25_ (.D(n1900),
	.CK(CLK),
	.Q(REGISTERS[793]));
   DFF_X1 REGISTERS_reg_7__24_ (.D(n1899),
	.CK(CLK),
	.Q(REGISTERS[792]));
   DFF_X1 REGISTERS_reg_7__23_ (.D(n1898),
	.CK(CLK),
	.Q(REGISTERS[791]));
   DFF_X1 REGISTERS_reg_7__22_ (.D(n1897),
	.CK(CLK),
	.Q(REGISTERS[790]));
   DFF_X1 REGISTERS_reg_7__21_ (.D(n1896),
	.CK(CLK),
	.Q(REGISTERS[789]));
   DFF_X1 REGISTERS_reg_7__20_ (.D(n1895),
	.CK(CLK),
	.Q(REGISTERS[788]));
   DFF_X1 REGISTERS_reg_7__19_ (.D(n1894),
	.CK(CLK),
	.Q(REGISTERS[787]));
   DFF_X1 REGISTERS_reg_7__18_ (.D(n1893),
	.CK(CLK),
	.Q(REGISTERS[786]));
   DFF_X1 REGISTERS_reg_7__17_ (.D(n1892),
	.CK(CLK),
	.Q(REGISTERS[785]));
   DFF_X1 REGISTERS_reg_7__16_ (.D(n1891),
	.CK(CLK),
	.Q(REGISTERS[784]));
   DFF_X1 REGISTERS_reg_7__15_ (.D(n1890),
	.CK(CLK),
	.Q(REGISTERS[783]));
   DFF_X1 REGISTERS_reg_7__14_ (.D(n1889),
	.CK(CLK),
	.Q(REGISTERS[782]));
   DFF_X1 REGISTERS_reg_7__13_ (.D(n1888),
	.CK(CLK),
	.Q(REGISTERS[781]));
   DFF_X1 REGISTERS_reg_7__12_ (.D(n1887),
	.CK(CLK),
	.Q(REGISTERS[780]));
   DFF_X1 REGISTERS_reg_7__11_ (.D(n1886),
	.CK(CLK),
	.Q(REGISTERS[779]));
   DFF_X1 REGISTERS_reg_7__10_ (.D(n1885),
	.CK(CLK),
	.Q(REGISTERS[778]));
   DFF_X1 REGISTERS_reg_7__9_ (.D(n1884),
	.CK(CLK),
	.Q(REGISTERS[777]));
   DFF_X1 REGISTERS_reg_7__8_ (.D(n1883),
	.CK(CLK),
	.Q(REGISTERS[776]));
   DFF_X1 REGISTERS_reg_7__7_ (.D(n1882),
	.CK(CLK),
	.Q(REGISTERS[775]));
   DFF_X1 REGISTERS_reg_7__6_ (.D(n1881),
	.CK(CLK),
	.Q(REGISTERS[774]));
   DFF_X1 REGISTERS_reg_7__5_ (.D(n1880),
	.CK(CLK),
	.Q(REGISTERS[773]));
   DFF_X1 REGISTERS_reg_7__4_ (.D(n1879),
	.CK(CLK),
	.Q(REGISTERS[772]));
   DFF_X1 REGISTERS_reg_7__3_ (.D(n1878),
	.CK(CLK),
	.Q(REGISTERS[771]));
   DFF_X1 REGISTERS_reg_7__2_ (.D(n1877),
	.CK(CLK),
	.Q(REGISTERS[770]));
   DFF_X1 REGISTERS_reg_7__1_ (.D(n1876),
	.CK(CLK),
	.Q(REGISTERS[769]));
   DFF_X1 REGISTERS_reg_7__0_ (.D(n1875),
	.CK(CLK),
	.Q(REGISTERS[768]));
   DFF_X1 REGISTERS_reg_8__31_ (.D(n1874),
	.CK(CLK),
	.Q(REGISTERS[767]));
   DFF_X1 REGISTERS_reg_8__30_ (.D(n1873),
	.CK(CLK),
	.Q(REGISTERS[766]));
   DFF_X1 REGISTERS_reg_8__29_ (.D(n1872),
	.CK(CLK),
	.Q(REGISTERS[765]));
   DFF_X1 REGISTERS_reg_8__28_ (.D(n1871),
	.CK(CLK),
	.Q(REGISTERS[764]));
   DFF_X1 REGISTERS_reg_8__27_ (.D(n1870),
	.CK(CLK),
	.Q(REGISTERS[763]));
   DFF_X1 REGISTERS_reg_8__26_ (.D(n1869),
	.CK(CLK),
	.Q(REGISTERS[762]));
   DFF_X1 REGISTERS_reg_8__25_ (.D(n1868),
	.CK(CLK),
	.Q(REGISTERS[761]));
   DFF_X1 REGISTERS_reg_8__24_ (.D(n1867),
	.CK(CLK),
	.Q(REGISTERS[760]));
   DFF_X1 REGISTERS_reg_8__23_ (.D(n1866),
	.CK(CLK),
	.Q(REGISTERS[759]));
   DFF_X1 REGISTERS_reg_8__22_ (.D(n1865),
	.CK(CLK),
	.Q(REGISTERS[758]));
   DFF_X1 REGISTERS_reg_8__21_ (.D(n1864),
	.CK(CLK),
	.Q(REGISTERS[757]));
   DFF_X1 REGISTERS_reg_8__20_ (.D(n1863),
	.CK(CLK),
	.Q(REGISTERS[756]));
   DFF_X1 REGISTERS_reg_8__19_ (.D(n1862),
	.CK(CLK),
	.Q(REGISTERS[755]));
   DFF_X1 REGISTERS_reg_8__18_ (.D(n1861),
	.CK(CLK),
	.Q(REGISTERS[754]));
   DFF_X1 REGISTERS_reg_8__17_ (.D(n1860),
	.CK(CLK),
	.Q(REGISTERS[753]));
   DFF_X1 REGISTERS_reg_8__16_ (.D(n1859),
	.CK(CLK),
	.Q(REGISTERS[752]));
   DFF_X1 REGISTERS_reg_8__15_ (.D(n1858),
	.CK(CLK),
	.Q(REGISTERS[751]));
   DFF_X1 REGISTERS_reg_8__14_ (.D(n1857),
	.CK(CLK),
	.Q(REGISTERS[750]));
   DFF_X1 REGISTERS_reg_8__13_ (.D(n1856),
	.CK(CLK),
	.Q(REGISTERS[749]));
   DFF_X1 REGISTERS_reg_8__12_ (.D(n1855),
	.CK(CLK),
	.Q(REGISTERS[748]));
   DFF_X1 REGISTERS_reg_8__11_ (.D(n1854),
	.CK(CLK),
	.Q(REGISTERS[747]));
   DFF_X1 REGISTERS_reg_8__10_ (.D(n1853),
	.CK(CLK),
	.Q(REGISTERS[746]));
   DFF_X1 REGISTERS_reg_8__9_ (.D(n1852),
	.CK(CLK),
	.Q(REGISTERS[745]));
   DFF_X1 REGISTERS_reg_8__8_ (.D(n1851),
	.CK(CLK),
	.Q(REGISTERS[744]));
   DFF_X1 REGISTERS_reg_8__7_ (.D(n1850),
	.CK(CLK),
	.Q(REGISTERS[743]));
   DFF_X1 REGISTERS_reg_8__6_ (.D(n1849),
	.CK(CLK),
	.Q(REGISTERS[742]));
   DFF_X1 REGISTERS_reg_8__5_ (.D(n1848),
	.CK(CLK),
	.Q(REGISTERS[741]));
   DFF_X1 REGISTERS_reg_8__4_ (.D(n1847),
	.CK(CLK),
	.Q(REGISTERS[740]));
   DFF_X1 REGISTERS_reg_8__3_ (.D(n1846),
	.CK(CLK),
	.Q(REGISTERS[739]));
   DFF_X1 REGISTERS_reg_8__2_ (.D(n1845),
	.CK(CLK),
	.Q(REGISTERS[738]));
   DFF_X1 REGISTERS_reg_8__1_ (.D(n1844),
	.CK(CLK),
	.Q(REGISTERS[737]));
   DFF_X1 REGISTERS_reg_8__0_ (.D(n1843),
	.CK(CLK),
	.Q(REGISTERS[736]));
   DFF_X1 REGISTERS_reg_9__31_ (.D(n1842),
	.CK(CLK),
	.Q(REGISTERS[735]));
   DFF_X1 REGISTERS_reg_9__30_ (.D(n1841),
	.CK(CLK),
	.Q(REGISTERS[734]));
   DFF_X1 REGISTERS_reg_9__29_ (.D(n1840),
	.CK(CLK),
	.Q(REGISTERS[733]));
   DFF_X1 REGISTERS_reg_9__28_ (.D(n1839),
	.CK(CLK),
	.Q(REGISTERS[732]));
   DFF_X1 REGISTERS_reg_9__27_ (.D(n1838),
	.CK(CLK),
	.Q(REGISTERS[731]));
   DFF_X1 REGISTERS_reg_9__26_ (.D(n1837),
	.CK(CLK),
	.Q(REGISTERS[730]));
   DFF_X1 REGISTERS_reg_9__25_ (.D(n1836),
	.CK(CLK),
	.Q(REGISTERS[729]));
   DFF_X1 REGISTERS_reg_9__24_ (.D(n1835),
	.CK(CLK),
	.Q(REGISTERS[728]));
   DFF_X1 REGISTERS_reg_9__23_ (.D(n1834),
	.CK(CLK),
	.Q(REGISTERS[727]));
   DFF_X1 REGISTERS_reg_9__22_ (.D(n1833),
	.CK(CLK),
	.Q(REGISTERS[726]));
   DFF_X1 REGISTERS_reg_9__21_ (.D(n1832),
	.CK(CLK),
	.Q(REGISTERS[725]));
   DFF_X1 REGISTERS_reg_9__20_ (.D(n1831),
	.CK(CLK),
	.Q(REGISTERS[724]));
   DFF_X1 REGISTERS_reg_9__19_ (.D(n1830),
	.CK(CLK),
	.Q(REGISTERS[723]));
   DFF_X1 REGISTERS_reg_9__18_ (.D(n1829),
	.CK(CLK),
	.Q(REGISTERS[722]));
   DFF_X1 REGISTERS_reg_9__17_ (.D(n1828),
	.CK(CLK),
	.Q(REGISTERS[721]));
   DFF_X1 REGISTERS_reg_9__16_ (.D(n1827),
	.CK(CLK),
	.Q(REGISTERS[720]));
   DFF_X1 REGISTERS_reg_9__15_ (.D(n1826),
	.CK(CLK),
	.Q(REGISTERS[719]));
   DFF_X1 REGISTERS_reg_9__14_ (.D(n1825),
	.CK(CLK),
	.Q(REGISTERS[718]));
   DFF_X1 REGISTERS_reg_9__13_ (.D(n1824),
	.CK(CLK),
	.Q(REGISTERS[717]));
   DFF_X1 REGISTERS_reg_9__12_ (.D(n1823),
	.CK(CLK),
	.Q(REGISTERS[716]));
   DFF_X1 REGISTERS_reg_9__11_ (.D(n1822),
	.CK(CLK),
	.Q(REGISTERS[715]));
   DFF_X1 REGISTERS_reg_9__10_ (.D(n1821),
	.CK(CLK),
	.Q(REGISTERS[714]));
   DFF_X1 REGISTERS_reg_9__9_ (.D(n1820),
	.CK(CLK),
	.Q(REGISTERS[713]));
   DFF_X1 REGISTERS_reg_9__8_ (.D(n1819),
	.CK(CLK),
	.Q(REGISTERS[712]));
   DFF_X1 REGISTERS_reg_9__7_ (.D(n1818),
	.CK(CLK),
	.Q(REGISTERS[711]));
   DFF_X1 REGISTERS_reg_9__6_ (.D(n1817),
	.CK(CLK),
	.Q(REGISTERS[710]));
   DFF_X1 REGISTERS_reg_9__5_ (.D(n1816),
	.CK(CLK),
	.Q(REGISTERS[709]));
   DFF_X1 REGISTERS_reg_9__4_ (.D(n1815),
	.CK(CLK),
	.Q(REGISTERS[708]));
   DFF_X1 REGISTERS_reg_9__3_ (.D(n1814),
	.CK(CLK),
	.Q(REGISTERS[707]));
   DFF_X1 REGISTERS_reg_9__2_ (.D(n1813),
	.CK(CLK),
	.Q(REGISTERS[706]));
   DFF_X1 REGISTERS_reg_9__1_ (.D(n1812),
	.CK(CLK),
	.Q(REGISTERS[705]));
   DFF_X1 REGISTERS_reg_9__0_ (.D(n1811),
	.CK(CLK),
	.Q(REGISTERS[704]));
   DFF_X1 REGISTERS_reg_10__31_ (.D(n1810),
	.CK(CLK),
	.Q(REGISTERS[703]));
   DFF_X1 REGISTERS_reg_10__30_ (.D(n1809),
	.CK(CLK),
	.Q(REGISTERS[702]));
   DFF_X1 REGISTERS_reg_10__29_ (.D(n1808),
	.CK(CLK),
	.Q(REGISTERS[701]));
   DFF_X1 REGISTERS_reg_10__28_ (.D(n1807),
	.CK(CLK),
	.Q(REGISTERS[700]));
   DFF_X1 REGISTERS_reg_10__27_ (.D(n1806),
	.CK(CLK),
	.Q(REGISTERS[699]));
   DFF_X1 REGISTERS_reg_10__26_ (.D(n1805),
	.CK(CLK),
	.Q(REGISTERS[698]));
   DFF_X1 REGISTERS_reg_10__25_ (.D(n1804),
	.CK(CLK),
	.Q(REGISTERS[697]));
   DFF_X1 REGISTERS_reg_10__24_ (.D(n1803),
	.CK(CLK),
	.Q(REGISTERS[696]));
   DFF_X1 REGISTERS_reg_10__23_ (.D(n1802),
	.CK(CLK),
	.Q(REGISTERS[695]));
   DFF_X1 REGISTERS_reg_10__22_ (.D(n1801),
	.CK(CLK),
	.Q(REGISTERS[694]));
   DFF_X1 REGISTERS_reg_10__21_ (.D(n1800),
	.CK(CLK),
	.Q(REGISTERS[693]));
   DFF_X1 REGISTERS_reg_10__20_ (.D(n1799),
	.CK(CLK),
	.Q(REGISTERS[692]));
   DFF_X1 REGISTERS_reg_10__19_ (.D(n1798),
	.CK(CLK),
	.Q(REGISTERS[691]));
   DFF_X1 REGISTERS_reg_10__18_ (.D(n1797),
	.CK(CLK),
	.Q(REGISTERS[690]));
   DFF_X1 REGISTERS_reg_10__17_ (.D(n1796),
	.CK(CLK),
	.Q(REGISTERS[689]));
   DFF_X1 REGISTERS_reg_10__16_ (.D(n1795),
	.CK(CLK),
	.Q(REGISTERS[688]));
   DFF_X1 REGISTERS_reg_10__15_ (.D(n1794),
	.CK(CLK),
	.Q(REGISTERS[687]));
   DFF_X1 REGISTERS_reg_10__14_ (.D(n1793),
	.CK(CLK),
	.Q(REGISTERS[686]));
   DFF_X1 REGISTERS_reg_10__13_ (.D(n1792),
	.CK(CLK),
	.Q(REGISTERS[685]));
   DFF_X1 REGISTERS_reg_10__12_ (.D(n1791),
	.CK(CLK),
	.Q(REGISTERS[684]));
   DFF_X1 REGISTERS_reg_10__11_ (.D(n1790),
	.CK(CLK),
	.Q(REGISTERS[683]));
   DFF_X1 REGISTERS_reg_10__10_ (.D(n1789),
	.CK(CLK),
	.Q(REGISTERS[682]));
   DFF_X1 REGISTERS_reg_10__9_ (.D(n1788),
	.CK(CLK),
	.Q(REGISTERS[681]));
   DFF_X1 REGISTERS_reg_10__8_ (.D(n1787),
	.CK(CLK),
	.Q(REGISTERS[680]));
   DFF_X1 REGISTERS_reg_10__7_ (.D(n1786),
	.CK(CLK),
	.Q(REGISTERS[679]));
   DFF_X1 REGISTERS_reg_10__6_ (.D(n1785),
	.CK(CLK),
	.Q(REGISTERS[678]));
   DFF_X1 REGISTERS_reg_10__5_ (.D(n1784),
	.CK(CLK),
	.Q(REGISTERS[677]));
   DFF_X1 REGISTERS_reg_10__4_ (.D(n1783),
	.CK(CLK),
	.Q(REGISTERS[676]));
   DFF_X1 REGISTERS_reg_10__3_ (.D(n1782),
	.CK(CLK),
	.Q(REGISTERS[675]));
   DFF_X1 REGISTERS_reg_10__2_ (.D(n1781),
	.CK(CLK),
	.Q(REGISTERS[674]));
   DFF_X1 REGISTERS_reg_10__1_ (.D(n1780),
	.CK(CLK),
	.Q(REGISTERS[673]));
   DFF_X1 REGISTERS_reg_10__0_ (.D(n1779),
	.CK(CLK),
	.Q(REGISTERS[672]));
   DFF_X1 REGISTERS_reg_11__31_ (.D(n1778),
	.CK(CLK),
	.Q(REGISTERS[671]));
   DFF_X1 REGISTERS_reg_11__30_ (.D(n1777),
	.CK(CLK),
	.Q(REGISTERS[670]));
   DFF_X1 REGISTERS_reg_11__29_ (.D(n1776),
	.CK(CLK),
	.Q(REGISTERS[669]));
   DFF_X1 REGISTERS_reg_11__28_ (.D(n1775),
	.CK(CLK),
	.Q(REGISTERS[668]));
   DFF_X1 REGISTERS_reg_11__27_ (.D(n1774),
	.CK(CLK),
	.Q(REGISTERS[667]));
   DFF_X1 REGISTERS_reg_11__26_ (.D(n1773),
	.CK(CLK),
	.Q(REGISTERS[666]));
   DFF_X1 REGISTERS_reg_11__25_ (.D(n1772),
	.CK(CLK),
	.Q(REGISTERS[665]));
   DFF_X1 REGISTERS_reg_11__24_ (.D(n1771),
	.CK(CLK),
	.Q(REGISTERS[664]));
   DFF_X1 REGISTERS_reg_11__23_ (.D(n1770),
	.CK(CLK),
	.Q(REGISTERS[663]));
   DFF_X1 REGISTERS_reg_11__22_ (.D(n1769),
	.CK(CLK),
	.Q(REGISTERS[662]));
   DFF_X1 REGISTERS_reg_11__21_ (.D(n1768),
	.CK(CLK),
	.Q(REGISTERS[661]));
   DFF_X1 REGISTERS_reg_11__20_ (.D(n1767),
	.CK(CLK),
	.Q(REGISTERS[660]));
   DFF_X1 REGISTERS_reg_11__19_ (.D(n1766),
	.CK(CLK),
	.Q(REGISTERS[659]));
   DFF_X1 REGISTERS_reg_11__18_ (.D(n1765),
	.CK(CLK),
	.Q(REGISTERS[658]));
   DFF_X1 REGISTERS_reg_11__17_ (.D(n1764),
	.CK(CLK),
	.Q(REGISTERS[657]));
   DFF_X1 REGISTERS_reg_11__16_ (.D(n1763),
	.CK(CLK),
	.Q(REGISTERS[656]));
   DFF_X1 REGISTERS_reg_11__15_ (.D(n1762),
	.CK(CLK),
	.Q(REGISTERS[655]));
   DFF_X1 REGISTERS_reg_11__14_ (.D(n1761),
	.CK(CLK),
	.Q(REGISTERS[654]));
   DFF_X1 REGISTERS_reg_11__13_ (.D(n1760),
	.CK(CLK),
	.Q(REGISTERS[653]));
   DFF_X1 REGISTERS_reg_11__12_ (.D(n1759),
	.CK(CLK),
	.Q(REGISTERS[652]));
   DFF_X1 REGISTERS_reg_11__11_ (.D(n1758),
	.CK(CLK),
	.Q(REGISTERS[651]));
   DFF_X1 REGISTERS_reg_11__10_ (.D(n1757),
	.CK(CLK),
	.Q(REGISTERS[650]));
   DFF_X1 REGISTERS_reg_11__9_ (.D(n1756),
	.CK(CLK),
	.Q(REGISTERS[649]));
   DFF_X1 REGISTERS_reg_11__8_ (.D(n1755),
	.CK(CLK),
	.Q(REGISTERS[648]));
   DFF_X1 REGISTERS_reg_11__7_ (.D(n1754),
	.CK(CLK),
	.Q(REGISTERS[647]));
   DFF_X1 REGISTERS_reg_11__6_ (.D(n1753),
	.CK(CLK),
	.Q(REGISTERS[646]));
   DFF_X1 REGISTERS_reg_11__5_ (.D(n1752),
	.CK(CLK),
	.Q(REGISTERS[645]));
   DFF_X1 REGISTERS_reg_11__4_ (.D(n1751),
	.CK(CLK),
	.Q(REGISTERS[644]));
   DFF_X1 REGISTERS_reg_11__3_ (.D(n1750),
	.CK(CLK),
	.Q(REGISTERS[643]));
   DFF_X1 REGISTERS_reg_11__2_ (.D(n1749),
	.CK(CLK),
	.Q(REGISTERS[642]));
   DFF_X1 REGISTERS_reg_11__1_ (.D(n1748),
	.CK(CLK),
	.Q(REGISTERS[641]));
   DFF_X1 REGISTERS_reg_11__0_ (.D(n1747),
	.CK(CLK),
	.Q(REGISTERS[640]));
   DFF_X1 REGISTERS_reg_12__31_ (.D(n1746),
	.CK(CLK),
	.Q(REGISTERS[639]));
   DFF_X1 REGISTERS_reg_12__30_ (.D(n1745),
	.CK(CLK),
	.Q(REGISTERS[638]));
   DFF_X1 REGISTERS_reg_12__29_ (.D(n1744),
	.CK(CLK),
	.Q(REGISTERS[637]));
   DFF_X1 REGISTERS_reg_12__28_ (.D(n1743),
	.CK(CLK),
	.Q(REGISTERS[636]));
   DFF_X1 REGISTERS_reg_12__27_ (.D(n1742),
	.CK(CLK),
	.Q(REGISTERS[635]));
   DFF_X1 REGISTERS_reg_12__26_ (.D(n1741),
	.CK(CLK),
	.Q(REGISTERS[634]));
   DFF_X1 REGISTERS_reg_12__25_ (.D(n1740),
	.CK(CLK),
	.Q(REGISTERS[633]));
   DFF_X1 REGISTERS_reg_12__24_ (.D(n1739),
	.CK(CLK),
	.Q(REGISTERS[632]));
   DFF_X1 REGISTERS_reg_12__23_ (.D(n1738),
	.CK(CLK),
	.Q(REGISTERS[631]));
   DFF_X1 REGISTERS_reg_12__22_ (.D(n1737),
	.CK(CLK),
	.Q(REGISTERS[630]));
   DFF_X1 REGISTERS_reg_12__21_ (.D(n1736),
	.CK(CLK),
	.Q(REGISTERS[629]));
   DFF_X1 REGISTERS_reg_12__20_ (.D(n1735),
	.CK(CLK),
	.Q(REGISTERS[628]));
   DFF_X1 REGISTERS_reg_12__19_ (.D(n1734),
	.CK(CLK),
	.Q(REGISTERS[627]));
   DFF_X1 REGISTERS_reg_12__18_ (.D(n1733),
	.CK(CLK),
	.Q(REGISTERS[626]));
   DFF_X1 REGISTERS_reg_12__17_ (.D(n1732),
	.CK(CLK),
	.Q(REGISTERS[625]));
   DFF_X1 REGISTERS_reg_12__16_ (.D(n1731),
	.CK(CLK),
	.Q(REGISTERS[624]));
   DFF_X1 REGISTERS_reg_12__15_ (.D(n1730),
	.CK(CLK),
	.Q(REGISTERS[623]));
   DFF_X1 REGISTERS_reg_12__14_ (.D(n1729),
	.CK(CLK),
	.Q(REGISTERS[622]));
   DFF_X1 REGISTERS_reg_12__13_ (.D(n1728),
	.CK(CLK),
	.Q(REGISTERS[621]));
   DFF_X1 REGISTERS_reg_12__12_ (.D(n1727),
	.CK(CLK),
	.Q(REGISTERS[620]));
   DFF_X1 REGISTERS_reg_12__11_ (.D(n1726),
	.CK(CLK),
	.Q(REGISTERS[619]));
   DFF_X1 REGISTERS_reg_12__10_ (.D(n1725),
	.CK(CLK),
	.Q(REGISTERS[618]));
   DFF_X1 REGISTERS_reg_12__9_ (.D(n1724),
	.CK(CLK),
	.Q(REGISTERS[617]));
   DFF_X1 REGISTERS_reg_12__8_ (.D(n1723),
	.CK(CLK),
	.Q(REGISTERS[616]));
   DFF_X1 REGISTERS_reg_12__7_ (.D(n1722),
	.CK(CLK),
	.Q(REGISTERS[615]));
   DFF_X1 REGISTERS_reg_12__6_ (.D(n1721),
	.CK(CLK),
	.Q(REGISTERS[614]));
   DFF_X1 REGISTERS_reg_12__5_ (.D(n1720),
	.CK(CLK),
	.Q(REGISTERS[613]));
   DFF_X1 REGISTERS_reg_12__4_ (.D(n1719),
	.CK(CLK),
	.Q(REGISTERS[612]));
   DFF_X1 REGISTERS_reg_12__3_ (.D(n1718),
	.CK(CLK),
	.Q(REGISTERS[611]));
   DFF_X1 REGISTERS_reg_12__2_ (.D(n1717),
	.CK(CLK),
	.Q(REGISTERS[610]));
   DFF_X1 REGISTERS_reg_12__1_ (.D(n1716),
	.CK(CLK),
	.Q(REGISTERS[609]));
   DFF_X1 REGISTERS_reg_12__0_ (.D(n1715),
	.CK(CLK),
	.Q(REGISTERS[608]));
   DFF_X1 REGISTERS_reg_13__31_ (.D(n1714),
	.CK(CLK),
	.Q(REGISTERS[607]));
   DFF_X1 REGISTERS_reg_13__30_ (.D(n1713),
	.CK(CLK),
	.Q(REGISTERS[606]));
   DFF_X1 REGISTERS_reg_13__29_ (.D(n1712),
	.CK(CLK),
	.Q(REGISTERS[605]));
   DFF_X1 REGISTERS_reg_13__28_ (.D(n1711),
	.CK(CLK),
	.Q(REGISTERS[604]));
   DFF_X1 REGISTERS_reg_13__27_ (.D(n1710),
	.CK(CLK),
	.Q(REGISTERS[603]));
   DFF_X1 REGISTERS_reg_13__26_ (.D(n1709),
	.CK(CLK),
	.Q(REGISTERS[602]));
   DFF_X1 REGISTERS_reg_13__25_ (.D(n1708),
	.CK(CLK),
	.Q(REGISTERS[601]));
   DFF_X1 REGISTERS_reg_13__24_ (.D(n1707),
	.CK(CLK),
	.Q(REGISTERS[600]));
   DFF_X1 REGISTERS_reg_13__23_ (.D(n1706),
	.CK(CLK),
	.Q(REGISTERS[599]));
   DFF_X1 REGISTERS_reg_13__22_ (.D(n1705),
	.CK(CLK),
	.Q(REGISTERS[598]));
   DFF_X1 REGISTERS_reg_13__21_ (.D(n1704),
	.CK(CLK),
	.Q(REGISTERS[597]));
   DFF_X1 REGISTERS_reg_13__20_ (.D(n1703),
	.CK(CLK),
	.Q(REGISTERS[596]));
   DFF_X1 REGISTERS_reg_13__19_ (.D(n1702),
	.CK(CLK),
	.Q(REGISTERS[595]));
   DFF_X1 REGISTERS_reg_13__18_ (.D(n1701),
	.CK(CLK),
	.Q(REGISTERS[594]));
   DFF_X1 REGISTERS_reg_13__17_ (.D(n1700),
	.CK(CLK),
	.Q(REGISTERS[593]));
   DFF_X1 REGISTERS_reg_13__16_ (.D(n1699),
	.CK(CLK),
	.Q(REGISTERS[592]));
   DFF_X1 REGISTERS_reg_13__15_ (.D(n1698),
	.CK(CLK),
	.Q(REGISTERS[591]));
   DFF_X1 REGISTERS_reg_13__14_ (.D(n1697),
	.CK(CLK),
	.Q(REGISTERS[590]));
   DFF_X1 REGISTERS_reg_13__13_ (.D(n1696),
	.CK(CLK),
	.Q(REGISTERS[589]));
   DFF_X1 REGISTERS_reg_13__12_ (.D(n1695),
	.CK(CLK),
	.Q(REGISTERS[588]));
   DFF_X1 REGISTERS_reg_13__11_ (.D(n1694),
	.CK(CLK),
	.Q(REGISTERS[587]));
   DFF_X1 REGISTERS_reg_13__10_ (.D(n1693),
	.CK(CLK),
	.Q(REGISTERS[586]));
   DFF_X1 REGISTERS_reg_13__9_ (.D(n1692),
	.CK(CLK),
	.Q(REGISTERS[585]));
   DFF_X1 REGISTERS_reg_13__8_ (.D(n1691),
	.CK(CLK),
	.Q(REGISTERS[584]));
   DFF_X1 REGISTERS_reg_13__7_ (.D(n1690),
	.CK(CLK),
	.Q(REGISTERS[583]));
   DFF_X1 REGISTERS_reg_13__6_ (.D(n1689),
	.CK(CLK),
	.Q(REGISTERS[582]));
   DFF_X1 REGISTERS_reg_13__5_ (.D(n1688),
	.CK(CLK),
	.Q(REGISTERS[581]));
   DFF_X1 REGISTERS_reg_13__4_ (.D(n1687),
	.CK(CLK),
	.Q(REGISTERS[580]));
   DFF_X1 REGISTERS_reg_13__3_ (.D(n1686),
	.CK(CLK),
	.Q(REGISTERS[579]));
   DFF_X1 REGISTERS_reg_13__2_ (.D(n1685),
	.CK(CLK),
	.Q(REGISTERS[578]));
   DFF_X1 REGISTERS_reg_13__1_ (.D(n1684),
	.CK(CLK),
	.Q(REGISTERS[577]));
   DFF_X1 REGISTERS_reg_13__0_ (.D(n1683),
	.CK(CLK),
	.Q(REGISTERS[576]));
   DFF_X1 REGISTERS_reg_14__31_ (.D(n1682),
	.CK(CLK),
	.Q(REGISTERS[575]));
   DFF_X1 REGISTERS_reg_14__30_ (.D(n1681),
	.CK(CLK),
	.Q(REGISTERS[574]));
   DFF_X1 REGISTERS_reg_14__29_ (.D(n1680),
	.CK(CLK),
	.Q(REGISTERS[573]));
   DFF_X1 REGISTERS_reg_14__28_ (.D(n1679),
	.CK(CLK),
	.Q(REGISTERS[572]));
   DFF_X1 REGISTERS_reg_14__27_ (.D(n1678),
	.CK(CLK),
	.Q(REGISTERS[571]));
   DFF_X1 REGISTERS_reg_14__26_ (.D(n1677),
	.CK(CLK),
	.Q(REGISTERS[570]));
   DFF_X1 REGISTERS_reg_14__25_ (.D(n1676),
	.CK(CLK),
	.Q(REGISTERS[569]));
   DFF_X1 REGISTERS_reg_14__24_ (.D(n1675),
	.CK(CLK),
	.Q(REGISTERS[568]));
   DFF_X1 REGISTERS_reg_14__23_ (.D(n1674),
	.CK(CLK),
	.Q(REGISTERS[567]));
   DFF_X1 REGISTERS_reg_14__22_ (.D(n1673),
	.CK(CLK),
	.Q(REGISTERS[566]));
   DFF_X1 REGISTERS_reg_14__21_ (.D(n1672),
	.CK(CLK),
	.Q(REGISTERS[565]));
   DFF_X1 REGISTERS_reg_14__20_ (.D(n1671),
	.CK(CLK),
	.Q(REGISTERS[564]));
   DFF_X1 REGISTERS_reg_14__19_ (.D(n1670),
	.CK(CLK),
	.Q(REGISTERS[563]));
   DFF_X1 REGISTERS_reg_14__18_ (.D(n1669),
	.CK(CLK),
	.Q(REGISTERS[562]));
   DFF_X1 REGISTERS_reg_14__17_ (.D(n1668),
	.CK(CLK),
	.Q(REGISTERS[561]));
   DFF_X1 REGISTERS_reg_14__16_ (.D(n1667),
	.CK(CLK),
	.Q(REGISTERS[560]));
   DFF_X1 REGISTERS_reg_14__15_ (.D(n1666),
	.CK(CLK),
	.Q(REGISTERS[559]));
   DFF_X1 REGISTERS_reg_14__14_ (.D(n1665),
	.CK(CLK),
	.Q(REGISTERS[558]));
   DFF_X1 REGISTERS_reg_14__13_ (.D(n1664),
	.CK(CLK),
	.Q(REGISTERS[557]));
   DFF_X1 REGISTERS_reg_14__12_ (.D(n1663),
	.CK(CLK),
	.Q(REGISTERS[556]));
   DFF_X1 REGISTERS_reg_14__11_ (.D(n1662),
	.CK(CLK),
	.Q(REGISTERS[555]));
   DFF_X1 REGISTERS_reg_14__10_ (.D(n1661),
	.CK(CLK),
	.Q(REGISTERS[554]));
   DFF_X1 REGISTERS_reg_14__9_ (.D(n1660),
	.CK(CLK),
	.Q(REGISTERS[553]));
   DFF_X1 REGISTERS_reg_14__8_ (.D(n1659),
	.CK(CLK),
	.Q(REGISTERS[552]));
   DFF_X1 REGISTERS_reg_14__7_ (.D(n1658),
	.CK(CLK),
	.Q(REGISTERS[551]));
   DFF_X1 REGISTERS_reg_14__6_ (.D(n1657),
	.CK(CLK),
	.Q(REGISTERS[550]));
   DFF_X1 REGISTERS_reg_14__5_ (.D(n1656),
	.CK(CLK),
	.Q(REGISTERS[549]));
   DFF_X1 REGISTERS_reg_14__4_ (.D(n1655),
	.CK(CLK),
	.Q(REGISTERS[548]));
   DFF_X1 REGISTERS_reg_14__3_ (.D(n1654),
	.CK(CLK),
	.Q(REGISTERS[547]));
   DFF_X1 REGISTERS_reg_14__2_ (.D(n1653),
	.CK(CLK),
	.Q(REGISTERS[546]));
   DFF_X1 REGISTERS_reg_14__1_ (.D(n1652),
	.CK(CLK),
	.Q(REGISTERS[545]));
   DFF_X1 REGISTERS_reg_14__0_ (.D(n1651),
	.CK(CLK),
	.Q(REGISTERS[544]));
   DFF_X1 REGISTERS_reg_15__31_ (.D(n1650),
	.CK(CLK),
	.Q(REGISTERS[543]));
   DFF_X1 REGISTERS_reg_15__30_ (.D(n1649),
	.CK(CLK),
	.Q(REGISTERS[542]));
   DFF_X1 REGISTERS_reg_15__29_ (.D(n1648),
	.CK(CLK),
	.Q(REGISTERS[541]));
   DFF_X1 REGISTERS_reg_15__28_ (.D(n1647),
	.CK(CLK),
	.Q(REGISTERS[540]));
   DFF_X1 REGISTERS_reg_15__27_ (.D(n1646),
	.CK(CLK),
	.Q(REGISTERS[539]));
   DFF_X1 REGISTERS_reg_15__26_ (.D(n1645),
	.CK(CLK),
	.Q(REGISTERS[538]));
   DFF_X1 REGISTERS_reg_15__25_ (.D(n1644),
	.CK(CLK),
	.Q(REGISTERS[537]));
   DFF_X1 REGISTERS_reg_15__24_ (.D(n1643),
	.CK(CLK),
	.Q(REGISTERS[536]));
   DFF_X1 REGISTERS_reg_15__23_ (.D(n1642),
	.CK(CLK),
	.Q(REGISTERS[535]));
   DFF_X1 REGISTERS_reg_15__22_ (.D(n1641),
	.CK(CLK),
	.Q(REGISTERS[534]));
   DFF_X1 REGISTERS_reg_15__21_ (.D(n1640),
	.CK(CLK),
	.Q(REGISTERS[533]));
   DFF_X1 REGISTERS_reg_15__20_ (.D(n1639),
	.CK(CLK),
	.Q(REGISTERS[532]));
   DFF_X1 REGISTERS_reg_15__19_ (.D(n1638),
	.CK(CLK),
	.Q(REGISTERS[531]));
   DFF_X1 REGISTERS_reg_15__18_ (.D(n1637),
	.CK(CLK),
	.Q(REGISTERS[530]));
   DFF_X1 REGISTERS_reg_15__17_ (.D(n1636),
	.CK(CLK),
	.Q(REGISTERS[529]));
   DFF_X1 REGISTERS_reg_15__16_ (.D(n1635),
	.CK(CLK),
	.Q(REGISTERS[528]));
   DFF_X1 REGISTERS_reg_15__15_ (.D(n1634),
	.CK(CLK),
	.Q(REGISTERS[527]));
   DFF_X1 REGISTERS_reg_15__14_ (.D(n1633),
	.CK(CLK),
	.Q(REGISTERS[526]));
   DFF_X1 REGISTERS_reg_15__13_ (.D(n1632),
	.CK(CLK),
	.Q(REGISTERS[525]));
   DFF_X1 REGISTERS_reg_15__12_ (.D(n1631),
	.CK(CLK),
	.Q(REGISTERS[524]));
   DFF_X1 REGISTERS_reg_15__11_ (.D(n1630),
	.CK(CLK),
	.Q(REGISTERS[523]));
   DFF_X1 REGISTERS_reg_15__10_ (.D(n1629),
	.CK(CLK),
	.Q(REGISTERS[522]));
   DFF_X1 REGISTERS_reg_15__9_ (.D(n1628),
	.CK(CLK),
	.Q(REGISTERS[521]));
   DFF_X1 REGISTERS_reg_15__8_ (.D(n1627),
	.CK(CLK),
	.Q(REGISTERS[520]));
   DFF_X1 REGISTERS_reg_15__7_ (.D(n1626),
	.CK(CLK),
	.Q(REGISTERS[519]));
   DFF_X1 REGISTERS_reg_15__6_ (.D(n1625),
	.CK(CLK),
	.Q(REGISTERS[518]));
   DFF_X1 REGISTERS_reg_15__5_ (.D(n1624),
	.CK(CLK),
	.Q(REGISTERS[517]));
   DFF_X1 REGISTERS_reg_15__4_ (.D(n1623),
	.CK(CLK),
	.Q(REGISTERS[516]));
   DFF_X1 REGISTERS_reg_15__3_ (.D(n1622),
	.CK(CLK),
	.Q(REGISTERS[515]));
   DFF_X1 REGISTERS_reg_15__2_ (.D(n1621),
	.CK(CLK),
	.Q(REGISTERS[514]));
   DFF_X1 REGISTERS_reg_15__1_ (.D(n1620),
	.CK(CLK),
	.Q(REGISTERS[513]));
   DFF_X1 REGISTERS_reg_15__0_ (.D(n1619),
	.CK(CLK),
	.Q(REGISTERS[512]));
   DFF_X1 REGISTERS_reg_16__31_ (.D(n1618),
	.CK(CLK),
	.Q(REGISTERS[511]));
   DFF_X1 REGISTERS_reg_16__30_ (.D(n1617),
	.CK(CLK),
	.Q(REGISTERS[510]));
   DFF_X1 REGISTERS_reg_16__29_ (.D(n1616),
	.CK(CLK),
	.Q(REGISTERS[509]));
   DFF_X1 REGISTERS_reg_16__28_ (.D(n1615),
	.CK(CLK),
	.Q(REGISTERS[508]));
   DFF_X1 REGISTERS_reg_16__27_ (.D(n1614),
	.CK(CLK),
	.Q(REGISTERS[507]));
   DFF_X1 REGISTERS_reg_16__26_ (.D(n1613),
	.CK(CLK),
	.Q(REGISTERS[506]));
   DFF_X1 REGISTERS_reg_16__25_ (.D(n1612),
	.CK(CLK),
	.Q(REGISTERS[505]));
   DFF_X1 REGISTERS_reg_16__24_ (.D(n1611),
	.CK(CLK),
	.Q(REGISTERS[504]));
   DFF_X1 REGISTERS_reg_16__23_ (.D(n1610),
	.CK(CLK),
	.Q(REGISTERS[503]));
   DFF_X1 REGISTERS_reg_16__22_ (.D(n1609),
	.CK(CLK),
	.Q(REGISTERS[502]));
   DFF_X1 REGISTERS_reg_16__21_ (.D(n1608),
	.CK(CLK),
	.Q(REGISTERS[501]));
   DFF_X1 REGISTERS_reg_16__20_ (.D(n1607),
	.CK(CLK),
	.Q(REGISTERS[500]));
   DFF_X1 REGISTERS_reg_16__19_ (.D(n1606),
	.CK(CLK),
	.Q(REGISTERS[499]));
   DFF_X1 REGISTERS_reg_16__18_ (.D(n1605),
	.CK(CLK),
	.Q(REGISTERS[498]));
   DFF_X1 REGISTERS_reg_16__17_ (.D(n1604),
	.CK(CLK),
	.Q(REGISTERS[497]));
   DFF_X1 REGISTERS_reg_16__16_ (.D(n1603),
	.CK(CLK),
	.Q(REGISTERS[496]));
   DFF_X1 REGISTERS_reg_16__15_ (.D(n1602),
	.CK(CLK),
	.Q(REGISTERS[495]));
   DFF_X1 REGISTERS_reg_16__14_ (.D(n1601),
	.CK(CLK),
	.Q(REGISTERS[494]));
   DFF_X1 REGISTERS_reg_16__13_ (.D(n1600),
	.CK(CLK),
	.Q(REGISTERS[493]));
   DFF_X1 REGISTERS_reg_16__12_ (.D(n1599),
	.CK(CLK),
	.Q(REGISTERS[492]));
   DFF_X1 REGISTERS_reg_16__11_ (.D(n1598),
	.CK(CLK),
	.Q(REGISTERS[491]));
   DFF_X1 REGISTERS_reg_16__10_ (.D(n1597),
	.CK(CLK),
	.Q(REGISTERS[490]));
   DFF_X1 REGISTERS_reg_16__9_ (.D(n1596),
	.CK(CLK),
	.Q(REGISTERS[489]));
   DFF_X1 REGISTERS_reg_16__8_ (.D(n1595),
	.CK(CLK),
	.Q(REGISTERS[488]));
   DFF_X1 REGISTERS_reg_16__7_ (.D(n1594),
	.CK(CLK),
	.Q(REGISTERS[487]));
   DFF_X1 REGISTERS_reg_16__6_ (.D(n1593),
	.CK(CLK),
	.Q(REGISTERS[486]));
   DFF_X1 REGISTERS_reg_16__5_ (.D(n1592),
	.CK(CLK),
	.Q(REGISTERS[485]));
   DFF_X1 REGISTERS_reg_16__4_ (.D(n1591),
	.CK(CLK),
	.Q(REGISTERS[484]));
   DFF_X1 REGISTERS_reg_16__3_ (.D(n1590),
	.CK(CLK),
	.Q(REGISTERS[483]));
   DFF_X1 REGISTERS_reg_16__2_ (.D(n1589),
	.CK(CLK),
	.Q(REGISTERS[482]));
   DFF_X1 REGISTERS_reg_16__1_ (.D(n1588),
	.CK(CLK),
	.Q(REGISTERS[481]));
   DFF_X1 REGISTERS_reg_16__0_ (.D(n1587),
	.CK(CLK),
	.Q(REGISTERS[480]));
   DFF_X1 REGISTERS_reg_17__31_ (.D(n1586),
	.CK(CLK),
	.Q(REGISTERS[479]));
   DFF_X1 REGISTERS_reg_17__30_ (.D(n1585),
	.CK(CLK),
	.Q(REGISTERS[478]));
   DFF_X1 REGISTERS_reg_17__29_ (.D(n1584),
	.CK(CLK),
	.Q(REGISTERS[477]));
   DFF_X1 REGISTERS_reg_17__28_ (.D(n1583),
	.CK(CLK),
	.Q(REGISTERS[476]));
   DFF_X1 REGISTERS_reg_17__27_ (.D(n1582),
	.CK(CLK),
	.Q(REGISTERS[475]));
   DFF_X1 REGISTERS_reg_17__26_ (.D(n1581),
	.CK(CLK),
	.Q(REGISTERS[474]));
   DFF_X1 REGISTERS_reg_17__25_ (.D(n1580),
	.CK(CLK),
	.Q(REGISTERS[473]));
   DFF_X1 REGISTERS_reg_17__24_ (.D(n1579),
	.CK(CLK),
	.Q(REGISTERS[472]));
   DFF_X1 REGISTERS_reg_17__23_ (.D(n1578),
	.CK(CLK),
	.Q(REGISTERS[471]));
   DFF_X1 REGISTERS_reg_17__22_ (.D(n1577),
	.CK(CLK),
	.Q(REGISTERS[470]));
   DFF_X1 REGISTERS_reg_17__21_ (.D(n1576),
	.CK(CLK),
	.Q(REGISTERS[469]));
   DFF_X1 REGISTERS_reg_17__20_ (.D(n1575),
	.CK(CLK),
	.Q(REGISTERS[468]));
   DFF_X1 REGISTERS_reg_17__19_ (.D(n1574),
	.CK(CLK),
	.Q(REGISTERS[467]));
   DFF_X1 REGISTERS_reg_17__18_ (.D(n1573),
	.CK(CLK),
	.Q(REGISTERS[466]));
   DFF_X1 REGISTERS_reg_17__17_ (.D(n1572),
	.CK(CLK),
	.Q(REGISTERS[465]));
   DFF_X1 REGISTERS_reg_17__16_ (.D(n1571),
	.CK(CLK),
	.Q(REGISTERS[464]));
   DFF_X1 REGISTERS_reg_17__15_ (.D(n1570),
	.CK(CLK),
	.Q(REGISTERS[463]));
   DFF_X1 REGISTERS_reg_17__14_ (.D(n1569),
	.CK(CLK),
	.Q(REGISTERS[462]));
   DFF_X1 REGISTERS_reg_17__13_ (.D(n1568),
	.CK(CLK),
	.Q(REGISTERS[461]));
   DFF_X1 REGISTERS_reg_17__12_ (.D(n1567),
	.CK(CLK),
	.Q(REGISTERS[460]));
   DFF_X1 REGISTERS_reg_17__11_ (.D(n1566),
	.CK(CLK),
	.Q(REGISTERS[459]));
   DFF_X1 REGISTERS_reg_17__10_ (.D(n1565),
	.CK(CLK),
	.Q(REGISTERS[458]));
   DFF_X1 REGISTERS_reg_17__9_ (.D(n1564),
	.CK(CLK),
	.Q(REGISTERS[457]));
   DFF_X1 REGISTERS_reg_17__8_ (.D(n1563),
	.CK(CLK),
	.Q(REGISTERS[456]));
   DFF_X1 REGISTERS_reg_17__7_ (.D(n1562),
	.CK(CLK),
	.Q(REGISTERS[455]));
   DFF_X1 REGISTERS_reg_17__6_ (.D(n1561),
	.CK(CLK),
	.Q(REGISTERS[454]));
   DFF_X1 REGISTERS_reg_17__5_ (.D(n1560),
	.CK(CLK),
	.Q(REGISTERS[453]));
   DFF_X1 REGISTERS_reg_17__4_ (.D(n1559),
	.CK(CLK),
	.Q(REGISTERS[452]));
   DFF_X1 REGISTERS_reg_17__3_ (.D(n1558),
	.CK(CLK),
	.Q(REGISTERS[451]));
   DFF_X1 REGISTERS_reg_17__2_ (.D(n1557),
	.CK(CLK),
	.Q(REGISTERS[450]));
   DFF_X1 REGISTERS_reg_17__1_ (.D(n1556),
	.CK(CLK),
	.Q(REGISTERS[449]));
   DFF_X1 REGISTERS_reg_17__0_ (.D(n1555),
	.CK(CLK),
	.Q(REGISTERS[448]));
   DFF_X1 REGISTERS_reg_18__31_ (.D(n1554),
	.CK(CLK),
	.Q(REGISTERS[447]));
   DFF_X1 REGISTERS_reg_18__30_ (.D(n1553),
	.CK(CLK),
	.Q(REGISTERS[446]));
   DFF_X1 REGISTERS_reg_18__29_ (.D(n1552),
	.CK(CLK),
	.Q(REGISTERS[445]));
   DFF_X1 REGISTERS_reg_18__28_ (.D(n1551),
	.CK(CLK),
	.Q(REGISTERS[444]));
   DFF_X1 REGISTERS_reg_18__27_ (.D(n1550),
	.CK(CLK),
	.Q(REGISTERS[443]));
   DFF_X1 REGISTERS_reg_18__26_ (.D(n1549),
	.CK(CLK),
	.Q(REGISTERS[442]));
   DFF_X1 REGISTERS_reg_18__25_ (.D(n1548),
	.CK(CLK),
	.Q(REGISTERS[441]));
   DFF_X1 REGISTERS_reg_18__24_ (.D(n1547),
	.CK(CLK),
	.Q(REGISTERS[440]));
   DFF_X1 REGISTERS_reg_18__23_ (.D(n1546),
	.CK(CLK),
	.Q(REGISTERS[439]));
   DFF_X1 REGISTERS_reg_18__22_ (.D(n1545),
	.CK(CLK),
	.Q(REGISTERS[438]));
   DFF_X1 REGISTERS_reg_18__21_ (.D(n1544),
	.CK(CLK),
	.Q(REGISTERS[437]));
   DFF_X1 REGISTERS_reg_18__20_ (.D(n1543),
	.CK(CLK),
	.Q(REGISTERS[436]));
   DFF_X1 REGISTERS_reg_18__19_ (.D(n1542),
	.CK(CLK),
	.Q(REGISTERS[435]));
   DFF_X1 REGISTERS_reg_18__18_ (.D(n1541),
	.CK(CLK),
	.Q(REGISTERS[434]));
   DFF_X1 REGISTERS_reg_18__17_ (.D(n1540),
	.CK(CLK),
	.Q(REGISTERS[433]));
   DFF_X1 REGISTERS_reg_18__16_ (.D(n1539),
	.CK(CLK),
	.Q(REGISTERS[432]));
   DFF_X1 REGISTERS_reg_18__15_ (.D(n1538),
	.CK(CLK),
	.Q(REGISTERS[431]));
   DFF_X1 REGISTERS_reg_18__14_ (.D(n1537),
	.CK(CLK),
	.Q(REGISTERS[430]));
   DFF_X1 REGISTERS_reg_18__13_ (.D(n1536),
	.CK(CLK),
	.Q(REGISTERS[429]));
   DFF_X1 REGISTERS_reg_18__12_ (.D(n1535),
	.CK(CLK),
	.Q(REGISTERS[428]));
   DFF_X1 REGISTERS_reg_18__11_ (.D(n1534),
	.CK(CLK),
	.Q(REGISTERS[427]));
   DFF_X1 REGISTERS_reg_18__10_ (.D(n1533),
	.CK(CLK),
	.Q(REGISTERS[426]));
   DFF_X1 REGISTERS_reg_18__9_ (.D(n1532),
	.CK(CLK),
	.Q(REGISTERS[425]));
   DFF_X1 REGISTERS_reg_18__8_ (.D(n1531),
	.CK(CLK),
	.Q(REGISTERS[424]));
   DFF_X1 REGISTERS_reg_18__7_ (.D(n1530),
	.CK(CLK),
	.Q(REGISTERS[423]));
   DFF_X1 REGISTERS_reg_18__6_ (.D(n1529),
	.CK(CLK),
	.Q(REGISTERS[422]));
   DFF_X1 REGISTERS_reg_18__5_ (.D(n1528),
	.CK(CLK),
	.Q(REGISTERS[421]));
   DFF_X1 REGISTERS_reg_18__4_ (.D(n1527),
	.CK(CLK),
	.Q(REGISTERS[420]));
   DFF_X1 REGISTERS_reg_18__3_ (.D(n1526),
	.CK(CLK),
	.Q(REGISTERS[419]));
   DFF_X1 REGISTERS_reg_18__2_ (.D(n1525),
	.CK(CLK),
	.Q(REGISTERS[418]));
   DFF_X1 REGISTERS_reg_18__1_ (.D(n1524),
	.CK(CLK),
	.Q(REGISTERS[417]));
   DFF_X1 REGISTERS_reg_18__0_ (.D(n1523),
	.CK(CLK),
	.Q(REGISTERS[416]));
   DFF_X1 REGISTERS_reg_19__31_ (.D(n1522),
	.CK(CLK),
	.Q(REGISTERS[415]));
   DFF_X1 REGISTERS_reg_19__30_ (.D(n1521),
	.CK(CLK),
	.Q(REGISTERS[414]));
   DFF_X1 REGISTERS_reg_19__29_ (.D(n1520),
	.CK(CLK),
	.Q(REGISTERS[413]));
   DFF_X1 REGISTERS_reg_19__28_ (.D(n1519),
	.CK(CLK),
	.Q(REGISTERS[412]));
   DFF_X1 REGISTERS_reg_19__27_ (.D(n1518),
	.CK(CLK),
	.Q(REGISTERS[411]));
   DFF_X1 REGISTERS_reg_19__26_ (.D(n1517),
	.CK(CLK),
	.Q(REGISTERS[410]));
   DFF_X1 REGISTERS_reg_19__25_ (.D(n1516),
	.CK(CLK),
	.Q(REGISTERS[409]));
   DFF_X1 REGISTERS_reg_19__24_ (.D(n1515),
	.CK(CLK),
	.Q(REGISTERS[408]));
   DFF_X1 REGISTERS_reg_19__23_ (.D(n1514),
	.CK(CLK),
	.Q(REGISTERS[407]));
   DFF_X1 REGISTERS_reg_19__22_ (.D(n1513),
	.CK(CLK),
	.Q(REGISTERS[406]));
   DFF_X1 REGISTERS_reg_19__21_ (.D(n1512),
	.CK(CLK),
	.Q(REGISTERS[405]));
   DFF_X1 REGISTERS_reg_19__20_ (.D(n1511),
	.CK(CLK),
	.Q(REGISTERS[404]));
   DFF_X1 REGISTERS_reg_19__19_ (.D(n1510),
	.CK(CLK),
	.Q(REGISTERS[403]));
   DFF_X1 REGISTERS_reg_19__18_ (.D(n1509),
	.CK(CLK),
	.Q(REGISTERS[402]));
   DFF_X1 REGISTERS_reg_19__17_ (.D(n1508),
	.CK(CLK),
	.Q(REGISTERS[401]));
   DFF_X1 REGISTERS_reg_19__16_ (.D(n1507),
	.CK(CLK),
	.Q(REGISTERS[400]));
   DFF_X1 REGISTERS_reg_19__15_ (.D(n1506),
	.CK(CLK),
	.Q(REGISTERS[399]));
   DFF_X1 REGISTERS_reg_19__14_ (.D(n1505),
	.CK(CLK),
	.Q(REGISTERS[398]));
   DFF_X1 REGISTERS_reg_19__13_ (.D(n1504),
	.CK(CLK),
	.Q(REGISTERS[397]));
   DFF_X1 REGISTERS_reg_19__12_ (.D(n1503),
	.CK(CLK),
	.Q(REGISTERS[396]));
   DFF_X1 REGISTERS_reg_19__11_ (.D(n1502),
	.CK(CLK),
	.Q(REGISTERS[395]));
   DFF_X1 REGISTERS_reg_19__10_ (.D(n1501),
	.CK(CLK),
	.Q(REGISTERS[394]));
   DFF_X1 REGISTERS_reg_19__9_ (.D(n1500),
	.CK(CLK),
	.Q(REGISTERS[393]));
   DFF_X1 REGISTERS_reg_19__8_ (.D(n1499),
	.CK(CLK),
	.Q(REGISTERS[392]));
   DFF_X1 REGISTERS_reg_19__7_ (.D(n1498),
	.CK(CLK),
	.Q(REGISTERS[391]));
   DFF_X1 REGISTERS_reg_19__6_ (.D(n1497),
	.CK(CLK),
	.Q(REGISTERS[390]));
   DFF_X1 REGISTERS_reg_19__5_ (.D(n1496),
	.CK(CLK),
	.Q(REGISTERS[389]));
   DFF_X1 REGISTERS_reg_19__4_ (.D(n1495),
	.CK(CLK),
	.Q(REGISTERS[388]));
   DFF_X1 REGISTERS_reg_19__3_ (.D(n1494),
	.CK(CLK),
	.Q(REGISTERS[387]));
   DFF_X1 REGISTERS_reg_19__2_ (.D(n1493),
	.CK(CLK),
	.Q(REGISTERS[386]));
   DFF_X1 REGISTERS_reg_19__1_ (.D(n1492),
	.CK(CLK),
	.Q(REGISTERS[385]));
   DFF_X1 REGISTERS_reg_19__0_ (.D(n1491),
	.CK(CLK),
	.Q(REGISTERS[384]));
   DFF_X1 REGISTERS_reg_20__31_ (.D(n1490),
	.CK(CLK),
	.Q(REGISTERS[383]));
   DFF_X1 REGISTERS_reg_20__30_ (.D(n1489),
	.CK(CLK),
	.Q(REGISTERS[382]));
   DFF_X1 REGISTERS_reg_20__29_ (.D(n1488),
	.CK(CLK),
	.Q(REGISTERS[381]));
   DFF_X1 REGISTERS_reg_20__28_ (.D(n1487),
	.CK(CLK),
	.Q(REGISTERS[380]));
   DFF_X1 REGISTERS_reg_20__27_ (.D(n1486),
	.CK(CLK),
	.Q(REGISTERS[379]));
   DFF_X1 REGISTERS_reg_20__26_ (.D(n1485),
	.CK(CLK),
	.Q(REGISTERS[378]));
   DFF_X1 REGISTERS_reg_20__25_ (.D(n1484),
	.CK(CLK),
	.Q(REGISTERS[377]));
   DFF_X1 REGISTERS_reg_20__24_ (.D(n1483),
	.CK(CLK),
	.Q(REGISTERS[376]));
   DFF_X1 REGISTERS_reg_20__23_ (.D(n1482),
	.CK(CLK),
	.Q(REGISTERS[375]));
   DFF_X1 REGISTERS_reg_20__22_ (.D(n1481),
	.CK(CLK),
	.Q(REGISTERS[374]));
   DFF_X1 REGISTERS_reg_20__21_ (.D(n1480),
	.CK(CLK),
	.Q(REGISTERS[373]));
   DFF_X1 REGISTERS_reg_20__20_ (.D(n1479),
	.CK(CLK),
	.Q(REGISTERS[372]));
   DFF_X1 REGISTERS_reg_20__19_ (.D(n1478),
	.CK(CLK),
	.Q(REGISTERS[371]));
   DFF_X1 REGISTERS_reg_20__18_ (.D(n1477),
	.CK(CLK),
	.Q(REGISTERS[370]));
   DFF_X1 REGISTERS_reg_20__17_ (.D(n1476),
	.CK(CLK),
	.Q(REGISTERS[369]));
   DFF_X1 REGISTERS_reg_20__16_ (.D(n1475),
	.CK(CLK),
	.Q(REGISTERS[368]));
   DFF_X1 REGISTERS_reg_20__15_ (.D(n1474),
	.CK(CLK),
	.Q(REGISTERS[367]));
   DFF_X1 REGISTERS_reg_20__14_ (.D(n1473),
	.CK(CLK),
	.Q(REGISTERS[366]));
   DFF_X1 REGISTERS_reg_20__13_ (.D(n1472),
	.CK(CLK),
	.Q(REGISTERS[365]));
   DFF_X1 REGISTERS_reg_20__12_ (.D(n1471),
	.CK(CLK),
	.Q(REGISTERS[364]));
   DFF_X1 REGISTERS_reg_20__11_ (.D(n1470),
	.CK(CLK),
	.Q(REGISTERS[363]));
   DFF_X1 REGISTERS_reg_20__10_ (.D(n1469),
	.CK(CLK),
	.Q(REGISTERS[362]));
   DFF_X1 REGISTERS_reg_20__9_ (.D(n1468),
	.CK(CLK),
	.Q(REGISTERS[361]));
   DFF_X1 REGISTERS_reg_20__8_ (.D(n1467),
	.CK(CLK),
	.Q(REGISTERS[360]));
   DFF_X1 REGISTERS_reg_20__7_ (.D(n1466),
	.CK(CLK),
	.Q(REGISTERS[359]));
   DFF_X1 REGISTERS_reg_20__6_ (.D(n1465),
	.CK(CLK),
	.Q(REGISTERS[358]));
   DFF_X1 REGISTERS_reg_20__5_ (.D(n1464),
	.CK(CLK),
	.Q(REGISTERS[357]));
   DFF_X1 REGISTERS_reg_20__4_ (.D(n1463),
	.CK(CLK),
	.Q(REGISTERS[356]));
   DFF_X1 REGISTERS_reg_20__3_ (.D(n1462),
	.CK(CLK),
	.Q(REGISTERS[355]));
   DFF_X1 REGISTERS_reg_20__2_ (.D(n1461),
	.CK(CLK),
	.Q(REGISTERS[354]));
   DFF_X1 REGISTERS_reg_20__1_ (.D(n1460),
	.CK(CLK),
	.Q(REGISTERS[353]));
   DFF_X1 REGISTERS_reg_20__0_ (.D(n1459),
	.CK(CLK),
	.Q(REGISTERS[352]));
   DFF_X1 REGISTERS_reg_21__31_ (.D(n1458),
	.CK(CLK),
	.Q(REGISTERS[351]));
   DFF_X1 REGISTERS_reg_21__30_ (.D(n1457),
	.CK(CLK),
	.Q(REGISTERS[350]));
   DFF_X1 REGISTERS_reg_21__29_ (.D(n1456),
	.CK(CLK),
	.Q(REGISTERS[349]));
   DFF_X1 REGISTERS_reg_21__28_ (.D(n1455),
	.CK(CLK),
	.Q(REGISTERS[348]));
   DFF_X1 REGISTERS_reg_21__27_ (.D(n1454),
	.CK(CLK),
	.Q(REGISTERS[347]));
   DFF_X1 REGISTERS_reg_21__26_ (.D(n1453),
	.CK(CLK),
	.Q(REGISTERS[346]));
   DFF_X1 REGISTERS_reg_21__25_ (.D(n1452),
	.CK(CLK),
	.Q(REGISTERS[345]));
   DFF_X1 REGISTERS_reg_21__24_ (.D(n1451),
	.CK(CLK),
	.Q(REGISTERS[344]));
   DFF_X1 REGISTERS_reg_21__23_ (.D(n1450),
	.CK(CLK),
	.Q(REGISTERS[343]));
   DFF_X1 REGISTERS_reg_21__22_ (.D(n1449),
	.CK(CLK),
	.Q(REGISTERS[342]));
   DFF_X1 REGISTERS_reg_21__21_ (.D(n1448),
	.CK(CLK),
	.Q(REGISTERS[341]));
   DFF_X1 REGISTERS_reg_21__20_ (.D(n1447),
	.CK(CLK),
	.Q(REGISTERS[340]));
   DFF_X1 REGISTERS_reg_21__19_ (.D(n1446),
	.CK(CLK),
	.Q(REGISTERS[339]));
   DFF_X1 REGISTERS_reg_21__18_ (.D(n1445),
	.CK(CLK),
	.Q(REGISTERS[338]));
   DFF_X1 REGISTERS_reg_21__17_ (.D(n1444),
	.CK(CLK),
	.Q(REGISTERS[337]));
   DFF_X1 REGISTERS_reg_21__16_ (.D(n1443),
	.CK(CLK),
	.Q(REGISTERS[336]));
   DFF_X1 REGISTERS_reg_21__15_ (.D(n1442),
	.CK(CLK),
	.Q(REGISTERS[335]));
   DFF_X1 REGISTERS_reg_21__14_ (.D(n1441),
	.CK(CLK),
	.Q(REGISTERS[334]));
   DFF_X1 REGISTERS_reg_21__13_ (.D(n1440),
	.CK(CLK),
	.Q(REGISTERS[333]));
   DFF_X1 REGISTERS_reg_21__12_ (.D(n1439),
	.CK(CLK),
	.Q(REGISTERS[332]));
   DFF_X1 REGISTERS_reg_21__11_ (.D(n1438),
	.CK(CLK),
	.Q(REGISTERS[331]));
   DFF_X1 REGISTERS_reg_21__10_ (.D(n1437),
	.CK(CLK),
	.Q(REGISTERS[330]));
   DFF_X1 REGISTERS_reg_21__9_ (.D(n1436),
	.CK(CLK),
	.Q(REGISTERS[329]));
   DFF_X1 REGISTERS_reg_21__8_ (.D(n1435),
	.CK(CLK),
	.Q(REGISTERS[328]));
   DFF_X1 REGISTERS_reg_21__7_ (.D(n1434),
	.CK(CLK),
	.Q(REGISTERS[327]));
   DFF_X1 REGISTERS_reg_21__6_ (.D(n1433),
	.CK(CLK),
	.Q(REGISTERS[326]));
   DFF_X1 REGISTERS_reg_21__5_ (.D(n1432),
	.CK(CLK),
	.Q(REGISTERS[325]));
   DFF_X1 REGISTERS_reg_21__4_ (.D(n1431),
	.CK(CLK),
	.Q(REGISTERS[324]));
   DFF_X1 REGISTERS_reg_21__3_ (.D(n1430),
	.CK(CLK),
	.Q(REGISTERS[323]));
   DFF_X1 REGISTERS_reg_21__2_ (.D(n1429),
	.CK(CLK),
	.Q(REGISTERS[322]));
   DFF_X1 REGISTERS_reg_21__1_ (.D(n1428),
	.CK(CLK),
	.Q(REGISTERS[321]));
   DFF_X1 REGISTERS_reg_21__0_ (.D(n1427),
	.CK(CLK),
	.Q(REGISTERS[320]));
   DFF_X1 REGISTERS_reg_22__31_ (.D(n1426),
	.CK(CLK),
	.Q(REGISTERS[319]));
   DFF_X1 REGISTERS_reg_22__30_ (.D(n1425),
	.CK(CLK),
	.Q(REGISTERS[318]));
   DFF_X1 REGISTERS_reg_22__29_ (.D(n1424),
	.CK(CLK),
	.Q(REGISTERS[317]));
   DFF_X1 REGISTERS_reg_22__28_ (.D(n1423),
	.CK(CLK),
	.Q(REGISTERS[316]));
   DFF_X1 REGISTERS_reg_22__27_ (.D(n1422),
	.CK(CLK),
	.Q(REGISTERS[315]));
   DFF_X1 REGISTERS_reg_22__26_ (.D(n1421),
	.CK(CLK),
	.Q(REGISTERS[314]));
   DFF_X1 REGISTERS_reg_22__25_ (.D(n1420),
	.CK(CLK),
	.Q(REGISTERS[313]));
   DFF_X1 REGISTERS_reg_22__24_ (.D(n1419),
	.CK(CLK),
	.Q(REGISTERS[312]));
   DFF_X1 REGISTERS_reg_22__23_ (.D(n1418),
	.CK(CLK),
	.Q(REGISTERS[311]));
   DFF_X1 REGISTERS_reg_22__22_ (.D(n1417),
	.CK(CLK),
	.Q(REGISTERS[310]));
   DFF_X1 REGISTERS_reg_22__21_ (.D(n1416),
	.CK(CLK),
	.Q(REGISTERS[309]));
   DFF_X1 REGISTERS_reg_22__20_ (.D(n1415),
	.CK(CLK),
	.Q(REGISTERS[308]));
   DFF_X1 REGISTERS_reg_22__19_ (.D(n1414),
	.CK(CLK),
	.Q(REGISTERS[307]));
   DFF_X1 REGISTERS_reg_22__18_ (.D(n1413),
	.CK(CLK),
	.Q(REGISTERS[306]));
   DFF_X1 REGISTERS_reg_22__17_ (.D(n1412),
	.CK(CLK),
	.Q(REGISTERS[305]));
   DFF_X1 REGISTERS_reg_22__16_ (.D(n1411),
	.CK(CLK),
	.Q(REGISTERS[304]));
   DFF_X1 REGISTERS_reg_22__15_ (.D(n1410),
	.CK(CLK),
	.Q(REGISTERS[303]));
   DFF_X1 REGISTERS_reg_22__14_ (.D(n1409),
	.CK(CLK),
	.Q(REGISTERS[302]));
   DFF_X1 REGISTERS_reg_22__13_ (.D(n1408),
	.CK(CLK),
	.Q(REGISTERS[301]));
   DFF_X1 REGISTERS_reg_22__12_ (.D(n1407),
	.CK(CLK),
	.Q(REGISTERS[300]));
   DFF_X1 REGISTERS_reg_22__11_ (.D(n1406),
	.CK(CLK),
	.Q(REGISTERS[299]));
   DFF_X1 REGISTERS_reg_22__10_ (.D(n1405),
	.CK(CLK),
	.Q(REGISTERS[298]));
   DFF_X1 REGISTERS_reg_22__9_ (.D(n1404),
	.CK(CLK),
	.Q(REGISTERS[297]));
   DFF_X1 REGISTERS_reg_22__8_ (.D(n1403),
	.CK(CLK),
	.Q(REGISTERS[296]));
   DFF_X1 REGISTERS_reg_22__7_ (.D(n1402),
	.CK(CLK),
	.Q(REGISTERS[295]));
   DFF_X1 REGISTERS_reg_22__6_ (.D(n1401),
	.CK(CLK),
	.Q(REGISTERS[294]));
   DFF_X1 REGISTERS_reg_22__5_ (.D(n1400),
	.CK(CLK),
	.Q(REGISTERS[293]));
   DFF_X1 REGISTERS_reg_22__4_ (.D(n1399),
	.CK(CLK),
	.Q(REGISTERS[292]));
   DFF_X1 REGISTERS_reg_22__3_ (.D(n1398),
	.CK(CLK),
	.Q(REGISTERS[291]));
   DFF_X1 REGISTERS_reg_22__2_ (.D(n1397),
	.CK(CLK),
	.Q(REGISTERS[290]));
   DFF_X1 REGISTERS_reg_22__1_ (.D(n1396),
	.CK(CLK),
	.Q(REGISTERS[289]));
   DFF_X1 REGISTERS_reg_22__0_ (.D(n1395),
	.CK(CLK),
	.Q(REGISTERS[288]));
   DFF_X1 REGISTERS_reg_23__31_ (.D(n1394),
	.CK(CLK),
	.Q(REGISTERS[287]));
   DFF_X1 REGISTERS_reg_23__30_ (.D(n1393),
	.CK(CLK),
	.Q(REGISTERS[286]));
   DFF_X1 REGISTERS_reg_23__29_ (.D(n1392),
	.CK(CLK),
	.Q(REGISTERS[285]));
   DFF_X1 REGISTERS_reg_23__28_ (.D(n1391),
	.CK(CLK),
	.Q(REGISTERS[284]));
   DFF_X1 REGISTERS_reg_23__27_ (.D(n1390),
	.CK(CLK),
	.Q(REGISTERS[283]));
   DFF_X1 REGISTERS_reg_23__26_ (.D(n1389),
	.CK(CLK),
	.Q(REGISTERS[282]));
   DFF_X1 REGISTERS_reg_23__25_ (.D(n1388),
	.CK(CLK),
	.Q(REGISTERS[281]));
   DFF_X1 REGISTERS_reg_23__24_ (.D(n1387),
	.CK(CLK),
	.Q(REGISTERS[280]));
   DFF_X1 REGISTERS_reg_23__23_ (.D(n1386),
	.CK(CLK),
	.Q(REGISTERS[279]));
   DFF_X1 REGISTERS_reg_23__22_ (.D(n1385),
	.CK(CLK),
	.Q(REGISTERS[278]));
   DFF_X1 REGISTERS_reg_23__21_ (.D(n1384),
	.CK(CLK),
	.Q(REGISTERS[277]));
   DFF_X1 REGISTERS_reg_23__20_ (.D(n1383),
	.CK(CLK),
	.Q(REGISTERS[276]));
   DFF_X1 REGISTERS_reg_23__19_ (.D(n1382),
	.CK(CLK),
	.Q(REGISTERS[275]));
   DFF_X1 REGISTERS_reg_23__18_ (.D(n1381),
	.CK(CLK),
	.Q(REGISTERS[274]));
   DFF_X1 REGISTERS_reg_23__17_ (.D(n1380),
	.CK(CLK),
	.Q(REGISTERS[273]));
   DFF_X1 REGISTERS_reg_23__16_ (.D(n1379),
	.CK(CLK),
	.Q(REGISTERS[272]));
   DFF_X1 REGISTERS_reg_23__15_ (.D(n1378),
	.CK(CLK),
	.Q(REGISTERS[271]));
   DFF_X1 REGISTERS_reg_23__14_ (.D(n1377),
	.CK(CLK),
	.Q(REGISTERS[270]));
   DFF_X1 REGISTERS_reg_23__13_ (.D(n1376),
	.CK(CLK),
	.Q(REGISTERS[269]));
   DFF_X1 REGISTERS_reg_23__12_ (.D(n1375),
	.CK(CLK),
	.Q(REGISTERS[268]));
   DFF_X1 REGISTERS_reg_23__11_ (.D(n1374),
	.CK(CLK),
	.Q(REGISTERS[267]));
   DFF_X1 REGISTERS_reg_23__10_ (.D(n1373),
	.CK(CLK),
	.Q(REGISTERS[266]));
   DFF_X1 REGISTERS_reg_23__9_ (.D(n1372),
	.CK(CLK),
	.Q(REGISTERS[265]));
   DFF_X1 REGISTERS_reg_23__8_ (.D(n1371),
	.CK(CLK),
	.Q(REGISTERS[264]));
   DFF_X1 REGISTERS_reg_23__7_ (.D(n1370),
	.CK(CLK),
	.Q(REGISTERS[263]));
   DFF_X1 REGISTERS_reg_23__6_ (.D(n1369),
	.CK(CLK),
	.Q(REGISTERS[262]));
   DFF_X1 REGISTERS_reg_23__5_ (.D(n1368),
	.CK(CLK),
	.Q(REGISTERS[261]));
   DFF_X1 REGISTERS_reg_23__4_ (.D(n1367),
	.CK(CLK),
	.Q(REGISTERS[260]));
   DFF_X1 REGISTERS_reg_23__3_ (.D(n1366),
	.CK(CLK),
	.Q(REGISTERS[259]));
   DFF_X1 REGISTERS_reg_23__2_ (.D(n1365),
	.CK(CLK),
	.Q(REGISTERS[258]));
   DFF_X1 REGISTERS_reg_23__1_ (.D(n1364),
	.CK(CLK),
	.Q(REGISTERS[257]));
   DFF_X1 REGISTERS_reg_23__0_ (.D(n1363),
	.CK(CLK),
	.Q(REGISTERS[256]));
   DFF_X1 REGISTERS_reg_24__31_ (.D(n1362),
	.CK(CLK),
	.Q(REGISTERS[255]));
   DFF_X1 REGISTERS_reg_24__30_ (.D(n1361),
	.CK(CLK),
	.Q(REGISTERS[254]));
   DFF_X1 REGISTERS_reg_24__29_ (.D(n1360),
	.CK(CLK),
	.Q(REGISTERS[253]));
   DFF_X1 REGISTERS_reg_24__28_ (.D(n1359),
	.CK(CLK),
	.Q(REGISTERS[252]));
   DFF_X1 REGISTERS_reg_24__27_ (.D(n1358),
	.CK(CLK),
	.Q(REGISTERS[251]));
   DFF_X1 REGISTERS_reg_24__26_ (.D(n1357),
	.CK(CLK),
	.Q(REGISTERS[250]));
   DFF_X1 REGISTERS_reg_24__25_ (.D(n1356),
	.CK(CLK),
	.Q(REGISTERS[249]));
   DFF_X1 REGISTERS_reg_24__24_ (.D(n1355),
	.CK(CLK),
	.Q(REGISTERS[248]));
   DFF_X1 REGISTERS_reg_24__23_ (.D(n1354),
	.CK(CLK),
	.Q(REGISTERS[247]));
   DFF_X1 REGISTERS_reg_24__22_ (.D(n1353),
	.CK(CLK),
	.Q(REGISTERS[246]));
   DFF_X1 REGISTERS_reg_24__21_ (.D(n1352),
	.CK(CLK),
	.Q(REGISTERS[245]));
   DFF_X1 REGISTERS_reg_24__20_ (.D(n1351),
	.CK(CLK),
	.Q(REGISTERS[244]));
   DFF_X1 REGISTERS_reg_24__19_ (.D(n1350),
	.CK(CLK),
	.Q(REGISTERS[243]));
   DFF_X1 REGISTERS_reg_24__18_ (.D(n1349),
	.CK(CLK),
	.Q(REGISTERS[242]));
   DFF_X1 REGISTERS_reg_24__17_ (.D(n1348),
	.CK(CLK),
	.Q(REGISTERS[241]));
   DFF_X1 REGISTERS_reg_24__16_ (.D(n1347),
	.CK(CLK),
	.Q(REGISTERS[240]));
   DFF_X1 REGISTERS_reg_24__15_ (.D(n1346),
	.CK(CLK),
	.Q(REGISTERS[239]));
   DFF_X1 REGISTERS_reg_24__14_ (.D(n1345),
	.CK(CLK),
	.Q(REGISTERS[238]));
   DFF_X1 REGISTERS_reg_24__13_ (.D(n1344),
	.CK(CLK),
	.Q(REGISTERS[237]));
   DFF_X1 REGISTERS_reg_24__12_ (.D(n1343),
	.CK(CLK),
	.Q(REGISTERS[236]));
   DFF_X1 REGISTERS_reg_24__11_ (.D(n1342),
	.CK(CLK),
	.Q(REGISTERS[235]));
   DFF_X1 REGISTERS_reg_24__10_ (.D(n1341),
	.CK(CLK),
	.Q(REGISTERS[234]));
   DFF_X1 REGISTERS_reg_24__9_ (.D(n1340),
	.CK(CLK),
	.Q(REGISTERS[233]));
   DFF_X1 REGISTERS_reg_24__8_ (.D(n1339),
	.CK(CLK),
	.Q(REGISTERS[232]));
   DFF_X1 REGISTERS_reg_24__7_ (.D(n1338),
	.CK(CLK),
	.Q(REGISTERS[231]));
   DFF_X1 REGISTERS_reg_24__6_ (.D(n1337),
	.CK(CLK),
	.Q(REGISTERS[230]));
   DFF_X1 REGISTERS_reg_24__5_ (.D(n1336),
	.CK(CLK),
	.Q(REGISTERS[229]));
   DFF_X1 REGISTERS_reg_24__4_ (.D(n1335),
	.CK(CLK),
	.Q(REGISTERS[228]));
   DFF_X1 REGISTERS_reg_24__3_ (.D(n1334),
	.CK(CLK),
	.Q(REGISTERS[227]));
   DFF_X1 REGISTERS_reg_24__2_ (.D(n1333),
	.CK(CLK),
	.Q(REGISTERS[226]));
   DFF_X1 REGISTERS_reg_24__1_ (.D(n1332),
	.CK(CLK),
	.Q(REGISTERS[225]));
   DFF_X1 REGISTERS_reg_24__0_ (.D(n1331),
	.CK(CLK),
	.Q(REGISTERS[224]));
   DFF_X1 REGISTERS_reg_25__31_ (.D(n1330),
	.CK(CLK),
	.Q(REGISTERS[223]));
   DFF_X1 REGISTERS_reg_25__30_ (.D(n1329),
	.CK(CLK),
	.Q(REGISTERS[222]));
   DFF_X1 REGISTERS_reg_25__29_ (.D(n1328),
	.CK(CLK),
	.Q(REGISTERS[221]));
   DFF_X1 REGISTERS_reg_25__28_ (.D(n1327),
	.CK(CLK),
	.Q(REGISTERS[220]));
   DFF_X1 REGISTERS_reg_25__27_ (.D(n1326),
	.CK(CLK),
	.Q(REGISTERS[219]));
   DFF_X1 REGISTERS_reg_25__26_ (.D(n1325),
	.CK(CLK),
	.Q(REGISTERS[218]));
   DFF_X1 REGISTERS_reg_25__25_ (.D(n1324),
	.CK(CLK),
	.Q(REGISTERS[217]));
   DFF_X1 REGISTERS_reg_25__24_ (.D(n1323),
	.CK(CLK),
	.Q(REGISTERS[216]));
   DFF_X1 REGISTERS_reg_25__23_ (.D(n1322),
	.CK(CLK),
	.Q(REGISTERS[215]));
   DFF_X1 REGISTERS_reg_25__22_ (.D(n1321),
	.CK(CLK),
	.Q(REGISTERS[214]));
   DFF_X1 REGISTERS_reg_25__21_ (.D(n1320),
	.CK(CLK),
	.Q(REGISTERS[213]));
   DFF_X1 REGISTERS_reg_25__20_ (.D(n1319),
	.CK(CLK),
	.Q(REGISTERS[212]));
   DFF_X1 REGISTERS_reg_25__19_ (.D(n1318),
	.CK(CLK),
	.Q(REGISTERS[211]));
   DFF_X1 REGISTERS_reg_25__18_ (.D(n1317),
	.CK(CLK),
	.Q(REGISTERS[210]));
   DFF_X1 REGISTERS_reg_25__17_ (.D(n1316),
	.CK(CLK),
	.Q(REGISTERS[209]));
   DFF_X1 REGISTERS_reg_25__16_ (.D(n1315),
	.CK(CLK),
	.Q(REGISTERS[208]));
   DFF_X1 REGISTERS_reg_25__15_ (.D(n1314),
	.CK(CLK),
	.Q(REGISTERS[207]));
   DFF_X1 REGISTERS_reg_25__14_ (.D(n1313),
	.CK(CLK),
	.Q(REGISTERS[206]));
   DFF_X1 REGISTERS_reg_25__13_ (.D(n1312),
	.CK(CLK),
	.Q(REGISTERS[205]));
   DFF_X1 REGISTERS_reg_25__12_ (.D(n1311),
	.CK(CLK),
	.Q(REGISTERS[204]));
   DFF_X1 REGISTERS_reg_25__11_ (.D(n1310),
	.CK(CLK),
	.Q(REGISTERS[203]));
   DFF_X1 REGISTERS_reg_25__10_ (.D(n1309),
	.CK(CLK),
	.Q(REGISTERS[202]));
   DFF_X1 REGISTERS_reg_25__9_ (.D(n1308),
	.CK(CLK),
	.Q(REGISTERS[201]));
   DFF_X1 REGISTERS_reg_25__8_ (.D(n1307),
	.CK(CLK),
	.Q(REGISTERS[200]));
   DFF_X1 REGISTERS_reg_25__7_ (.D(n1306),
	.CK(CLK),
	.Q(REGISTERS[199]));
   DFF_X1 REGISTERS_reg_25__6_ (.D(n1305),
	.CK(CLK),
	.Q(REGISTERS[198]));
   DFF_X1 REGISTERS_reg_25__5_ (.D(n1304),
	.CK(CLK),
	.Q(REGISTERS[197]));
   DFF_X1 REGISTERS_reg_25__4_ (.D(n1303),
	.CK(CLK),
	.Q(REGISTERS[196]));
   DFF_X1 REGISTERS_reg_25__3_ (.D(n1302),
	.CK(CLK),
	.Q(REGISTERS[195]));
   DFF_X1 REGISTERS_reg_25__2_ (.D(n1301),
	.CK(CLK),
	.Q(REGISTERS[194]));
   DFF_X1 REGISTERS_reg_25__1_ (.D(n1300),
	.CK(CLK),
	.Q(REGISTERS[193]));
   DFF_X1 REGISTERS_reg_25__0_ (.D(n1299),
	.CK(CLK),
	.Q(REGISTERS[192]));
   DFF_X1 REGISTERS_reg_26__31_ (.D(n1298),
	.CK(CLK),
	.Q(REGISTERS[191]));
   DFF_X1 REGISTERS_reg_26__30_ (.D(n1297),
	.CK(CLK),
	.Q(REGISTERS[190]));
   DFF_X1 REGISTERS_reg_26__29_ (.D(n1296),
	.CK(CLK),
	.Q(REGISTERS[189]));
   DFF_X1 REGISTERS_reg_26__28_ (.D(n1295),
	.CK(CLK),
	.Q(REGISTERS[188]));
   DFF_X1 REGISTERS_reg_26__27_ (.D(n1294),
	.CK(CLK),
	.Q(REGISTERS[187]));
   DFF_X1 REGISTERS_reg_26__26_ (.D(n1293),
	.CK(CLK),
	.Q(REGISTERS[186]));
   DFF_X1 REGISTERS_reg_26__25_ (.D(n1292),
	.CK(CLK),
	.Q(REGISTERS[185]));
   DFF_X1 REGISTERS_reg_26__24_ (.D(n1291),
	.CK(CLK),
	.Q(REGISTERS[184]));
   DFF_X1 REGISTERS_reg_26__23_ (.D(n1290),
	.CK(CLK),
	.Q(REGISTERS[183]));
   DFF_X1 REGISTERS_reg_26__22_ (.D(n1289),
	.CK(CLK),
	.Q(REGISTERS[182]));
   DFF_X1 REGISTERS_reg_26__21_ (.D(n1288),
	.CK(CLK),
	.Q(REGISTERS[181]));
   DFF_X1 REGISTERS_reg_26__20_ (.D(n1287),
	.CK(CLK),
	.Q(REGISTERS[180]));
   DFF_X1 REGISTERS_reg_26__19_ (.D(n1286),
	.CK(CLK),
	.Q(REGISTERS[179]));
   DFF_X1 REGISTERS_reg_26__18_ (.D(n1285),
	.CK(CLK),
	.Q(REGISTERS[178]));
   DFF_X1 REGISTERS_reg_26__17_ (.D(n1284),
	.CK(CLK),
	.Q(REGISTERS[177]));
   DFF_X1 REGISTERS_reg_26__16_ (.D(n1283),
	.CK(CLK),
	.Q(REGISTERS[176]));
   DFF_X1 REGISTERS_reg_26__15_ (.D(n1282),
	.CK(CLK),
	.Q(REGISTERS[175]));
   DFF_X1 REGISTERS_reg_26__14_ (.D(n1281),
	.CK(CLK),
	.Q(REGISTERS[174]));
   DFF_X1 REGISTERS_reg_26__13_ (.D(n1280),
	.CK(CLK),
	.Q(REGISTERS[173]));
   DFF_X1 REGISTERS_reg_26__12_ (.D(n1279),
	.CK(CLK),
	.Q(REGISTERS[172]));
   DFF_X1 REGISTERS_reg_26__11_ (.D(n1278),
	.CK(CLK),
	.Q(REGISTERS[171]));
   DFF_X1 REGISTERS_reg_26__10_ (.D(n1277),
	.CK(CLK),
	.Q(REGISTERS[170]));
   DFF_X1 REGISTERS_reg_26__9_ (.D(n1276),
	.CK(CLK),
	.Q(REGISTERS[169]));
   DFF_X1 REGISTERS_reg_26__8_ (.D(n1275),
	.CK(CLK),
	.Q(REGISTERS[168]));
   DFF_X1 REGISTERS_reg_26__7_ (.D(n1274),
	.CK(CLK),
	.Q(REGISTERS[167]));
   DFF_X1 REGISTERS_reg_26__6_ (.D(n1273),
	.CK(CLK),
	.Q(REGISTERS[166]));
   DFF_X1 REGISTERS_reg_26__5_ (.D(n1272),
	.CK(CLK),
	.Q(REGISTERS[165]));
   DFF_X1 REGISTERS_reg_26__4_ (.D(n1271),
	.CK(CLK),
	.Q(REGISTERS[164]));
   DFF_X1 REGISTERS_reg_26__3_ (.D(n1270),
	.CK(CLK),
	.Q(REGISTERS[163]));
   DFF_X1 REGISTERS_reg_26__2_ (.D(n1269),
	.CK(CLK),
	.Q(REGISTERS[162]));
   DFF_X1 REGISTERS_reg_26__1_ (.D(n1268),
	.CK(CLK),
	.Q(REGISTERS[161]));
   DFF_X1 REGISTERS_reg_26__0_ (.D(n1267),
	.CK(CLK),
	.Q(REGISTERS[160]));
   DFF_X1 REGISTERS_reg_27__31_ (.D(n1266),
	.CK(CLK),
	.Q(REGISTERS[159]));
   DFF_X1 REGISTERS_reg_27__30_ (.D(n1265),
	.CK(CLK),
	.Q(REGISTERS[158]));
   DFF_X1 REGISTERS_reg_27__29_ (.D(n1264),
	.CK(CLK),
	.Q(REGISTERS[157]));
   DFF_X1 REGISTERS_reg_27__28_ (.D(n1263),
	.CK(CLK),
	.Q(REGISTERS[156]));
   DFF_X1 REGISTERS_reg_27__27_ (.D(n1262),
	.CK(CLK),
	.Q(REGISTERS[155]));
   DFF_X1 REGISTERS_reg_27__26_ (.D(n1261),
	.CK(CLK),
	.Q(REGISTERS[154]));
   DFF_X1 REGISTERS_reg_27__25_ (.D(n1260),
	.CK(CLK),
	.Q(REGISTERS[153]));
   DFF_X1 REGISTERS_reg_27__24_ (.D(n1259),
	.CK(CLK),
	.Q(REGISTERS[152]));
   DFF_X1 REGISTERS_reg_27__23_ (.D(n1258),
	.CK(CLK),
	.Q(REGISTERS[151]));
   DFF_X1 REGISTERS_reg_27__22_ (.D(n1257),
	.CK(CLK),
	.Q(REGISTERS[150]));
   DFF_X1 REGISTERS_reg_27__21_ (.D(n1256),
	.CK(CLK),
	.Q(REGISTERS[149]));
   DFF_X1 REGISTERS_reg_27__20_ (.D(n1255),
	.CK(CLK),
	.Q(REGISTERS[148]));
   DFF_X1 REGISTERS_reg_27__19_ (.D(n1254),
	.CK(CLK),
	.Q(REGISTERS[147]));
   DFF_X1 REGISTERS_reg_27__18_ (.D(n1253),
	.CK(CLK),
	.Q(REGISTERS[146]));
   DFF_X1 REGISTERS_reg_27__17_ (.D(n1252),
	.CK(CLK),
	.Q(REGISTERS[145]));
   DFF_X1 REGISTERS_reg_27__16_ (.D(n1251),
	.CK(CLK),
	.Q(REGISTERS[144]));
   DFF_X1 REGISTERS_reg_27__15_ (.D(n1250),
	.CK(CLK),
	.Q(REGISTERS[143]));
   DFF_X1 REGISTERS_reg_27__14_ (.D(n1249),
	.CK(CLK),
	.Q(REGISTERS[142]));
   DFF_X1 REGISTERS_reg_27__13_ (.D(n1248),
	.CK(CLK),
	.Q(REGISTERS[141]));
   DFF_X1 REGISTERS_reg_27__12_ (.D(n1247),
	.CK(CLK),
	.Q(REGISTERS[140]));
   DFF_X1 REGISTERS_reg_27__11_ (.D(n1246),
	.CK(CLK),
	.Q(REGISTERS[139]));
   DFF_X1 REGISTERS_reg_27__10_ (.D(n1245),
	.CK(CLK),
	.Q(REGISTERS[138]));
   DFF_X1 REGISTERS_reg_27__9_ (.D(n1244),
	.CK(CLK),
	.Q(REGISTERS[137]));
   DFF_X1 REGISTERS_reg_27__8_ (.D(n1243),
	.CK(CLK),
	.Q(REGISTERS[136]));
   DFF_X1 REGISTERS_reg_27__7_ (.D(n1242),
	.CK(CLK),
	.Q(REGISTERS[135]));
   DFF_X1 REGISTERS_reg_27__6_ (.D(n1241),
	.CK(CLK),
	.Q(REGISTERS[134]));
   DFF_X1 REGISTERS_reg_27__5_ (.D(n1240),
	.CK(CLK),
	.Q(REGISTERS[133]));
   DFF_X1 REGISTERS_reg_27__4_ (.D(n1239),
	.CK(CLK),
	.Q(REGISTERS[132]));
   DFF_X1 REGISTERS_reg_27__3_ (.D(n1238),
	.CK(CLK),
	.Q(REGISTERS[131]));
   DFF_X1 REGISTERS_reg_27__2_ (.D(n1237),
	.CK(CLK),
	.Q(REGISTERS[130]));
   DFF_X1 REGISTERS_reg_27__1_ (.D(n1236),
	.CK(CLK),
	.Q(REGISTERS[129]));
   DFF_X1 REGISTERS_reg_27__0_ (.D(n1235),
	.CK(CLK),
	.Q(REGISTERS[128]));
   DFF_X1 REGISTERS_reg_28__31_ (.D(n1234),
	.CK(CLK),
	.Q(REGISTERS[127]));
   DFF_X1 REGISTERS_reg_28__30_ (.D(n1233),
	.CK(CLK),
	.Q(REGISTERS[126]));
   DFF_X1 REGISTERS_reg_28__29_ (.D(n1232),
	.CK(CLK),
	.Q(REGISTERS[125]));
   DFF_X1 REGISTERS_reg_28__28_ (.D(n1231),
	.CK(CLK),
	.Q(REGISTERS[124]));
   DFF_X1 REGISTERS_reg_28__27_ (.D(n1230),
	.CK(CLK),
	.Q(REGISTERS[123]));
   DFF_X1 REGISTERS_reg_28__26_ (.D(n1229),
	.CK(CLK),
	.Q(REGISTERS[122]));
   DFF_X1 REGISTERS_reg_28__25_ (.D(n1228),
	.CK(CLK),
	.Q(REGISTERS[121]));
   DFF_X1 REGISTERS_reg_28__24_ (.D(n1227),
	.CK(CLK),
	.Q(REGISTERS[120]));
   DFF_X1 REGISTERS_reg_28__23_ (.D(n1226),
	.CK(CLK),
	.Q(REGISTERS[119]));
   DFF_X1 REGISTERS_reg_28__22_ (.D(n1225),
	.CK(CLK),
	.Q(REGISTERS[118]));
   DFF_X1 REGISTERS_reg_28__21_ (.D(n1224),
	.CK(CLK),
	.Q(REGISTERS[117]));
   DFF_X1 REGISTERS_reg_28__20_ (.D(n1223),
	.CK(CLK),
	.Q(REGISTERS[116]));
   DFF_X1 REGISTERS_reg_28__19_ (.D(n1222),
	.CK(CLK),
	.Q(REGISTERS[115]));
   DFF_X1 REGISTERS_reg_28__18_ (.D(n1221),
	.CK(CLK),
	.Q(REGISTERS[114]));
   DFF_X1 REGISTERS_reg_28__17_ (.D(n1220),
	.CK(CLK),
	.Q(REGISTERS[113]));
   DFF_X1 REGISTERS_reg_28__16_ (.D(n1219),
	.CK(CLK),
	.Q(REGISTERS[112]));
   DFF_X1 REGISTERS_reg_28__15_ (.D(n1218),
	.CK(CLK),
	.Q(REGISTERS[111]));
   DFF_X1 REGISTERS_reg_28__14_ (.D(n1217),
	.CK(CLK),
	.Q(REGISTERS[110]));
   DFF_X1 REGISTERS_reg_28__13_ (.D(n1216),
	.CK(CLK),
	.Q(REGISTERS[109]));
   DFF_X1 REGISTERS_reg_28__12_ (.D(n1215),
	.CK(CLK),
	.Q(REGISTERS[108]));
   DFF_X1 REGISTERS_reg_28__11_ (.D(n1214),
	.CK(CLK),
	.Q(REGISTERS[107]));
   DFF_X1 REGISTERS_reg_28__10_ (.D(n1213),
	.CK(CLK),
	.Q(REGISTERS[106]));
   DFF_X1 REGISTERS_reg_28__9_ (.D(n1212),
	.CK(CLK),
	.Q(REGISTERS[105]));
   DFF_X1 REGISTERS_reg_28__8_ (.D(n1211),
	.CK(CLK),
	.Q(REGISTERS[104]));
   DFF_X1 REGISTERS_reg_28__7_ (.D(n1210),
	.CK(CLK),
	.Q(REGISTERS[103]));
   DFF_X1 REGISTERS_reg_28__6_ (.D(n1209),
	.CK(CLK),
	.Q(REGISTERS[102]));
   DFF_X1 REGISTERS_reg_28__5_ (.D(n1208),
	.CK(CLK),
	.Q(REGISTERS[101]));
   DFF_X1 REGISTERS_reg_28__4_ (.D(n1207),
	.CK(CLK),
	.Q(REGISTERS[100]));
   DFF_X1 REGISTERS_reg_28__3_ (.D(n1206),
	.CK(CLK),
	.Q(REGISTERS[99]));
   DFF_X1 REGISTERS_reg_28__2_ (.D(n1205),
	.CK(CLK),
	.Q(REGISTERS[98]));
   DFF_X1 REGISTERS_reg_28__1_ (.D(n1204),
	.CK(CLK),
	.Q(REGISTERS[97]));
   DFF_X1 REGISTERS_reg_28__0_ (.D(n1203),
	.CK(CLK),
	.Q(REGISTERS[96]));
   DFF_X1 REGISTERS_reg_29__31_ (.D(n1202),
	.CK(CLK),
	.Q(REGISTERS[95]));
   DFF_X1 REGISTERS_reg_29__30_ (.D(n1201),
	.CK(CLK),
	.Q(REGISTERS[94]));
   DFF_X1 REGISTERS_reg_29__29_ (.D(n1200),
	.CK(CLK),
	.Q(REGISTERS[93]));
   DFF_X1 REGISTERS_reg_29__28_ (.D(n1199),
	.CK(CLK),
	.Q(REGISTERS[92]));
   DFF_X1 REGISTERS_reg_29__27_ (.D(n1198),
	.CK(CLK),
	.Q(REGISTERS[91]));
   DFF_X1 REGISTERS_reg_29__26_ (.D(n1197),
	.CK(CLK),
	.Q(REGISTERS[90]));
   DFF_X1 REGISTERS_reg_29__25_ (.D(n1196),
	.CK(CLK),
	.Q(REGISTERS[89]));
   DFF_X1 REGISTERS_reg_29__24_ (.D(n1195),
	.CK(CLK),
	.Q(REGISTERS[88]));
   DFF_X1 REGISTERS_reg_29__23_ (.D(n1194),
	.CK(CLK),
	.Q(REGISTERS[87]));
   DFF_X1 REGISTERS_reg_29__22_ (.D(n1193),
	.CK(CLK),
	.Q(REGISTERS[86]));
   DFF_X1 REGISTERS_reg_29__21_ (.D(n1192),
	.CK(CLK),
	.Q(REGISTERS[85]));
   DFF_X1 REGISTERS_reg_29__20_ (.D(n1191),
	.CK(CLK),
	.Q(REGISTERS[84]));
   DFF_X1 REGISTERS_reg_29__19_ (.D(n1190),
	.CK(CLK),
	.Q(REGISTERS[83]));
   DFF_X1 REGISTERS_reg_29__18_ (.D(n1189),
	.CK(CLK),
	.Q(REGISTERS[82]));
   DFF_X1 REGISTERS_reg_29__17_ (.D(n1188),
	.CK(CLK),
	.Q(REGISTERS[81]));
   DFF_X1 REGISTERS_reg_29__16_ (.D(n1187),
	.CK(CLK),
	.Q(REGISTERS[80]));
   DFF_X1 REGISTERS_reg_29__15_ (.D(n1186),
	.CK(CLK),
	.Q(REGISTERS[79]));
   DFF_X1 REGISTERS_reg_29__14_ (.D(n1185),
	.CK(CLK),
	.Q(REGISTERS[78]));
   DFF_X1 REGISTERS_reg_29__13_ (.D(n1184),
	.CK(CLK),
	.Q(REGISTERS[77]));
   DFF_X1 REGISTERS_reg_29__12_ (.D(n1183),
	.CK(CLK),
	.Q(REGISTERS[76]));
   DFF_X1 REGISTERS_reg_29__11_ (.D(n1182),
	.CK(CLK),
	.Q(REGISTERS[75]));
   DFF_X1 REGISTERS_reg_29__10_ (.D(n1181),
	.CK(CLK),
	.Q(REGISTERS[74]));
   DFF_X1 REGISTERS_reg_29__9_ (.D(n1180),
	.CK(CLK),
	.Q(REGISTERS[73]));
   DFF_X1 REGISTERS_reg_29__8_ (.D(n1179),
	.CK(CLK),
	.Q(REGISTERS[72]));
   DFF_X1 REGISTERS_reg_29__7_ (.D(n1178),
	.CK(CLK),
	.Q(REGISTERS[71]));
   DFF_X1 REGISTERS_reg_29__6_ (.D(n1177),
	.CK(CLK),
	.Q(REGISTERS[70]));
   DFF_X1 REGISTERS_reg_29__5_ (.D(n1176),
	.CK(CLK),
	.Q(REGISTERS[69]));
   DFF_X1 REGISTERS_reg_29__4_ (.D(n1175),
	.CK(CLK),
	.Q(REGISTERS[68]));
   DFF_X1 REGISTERS_reg_29__3_ (.D(n1174),
	.CK(CLK),
	.Q(REGISTERS[67]));
   DFF_X1 REGISTERS_reg_29__2_ (.D(n1173),
	.CK(CLK),
	.Q(REGISTERS[66]));
   DFF_X1 REGISTERS_reg_29__1_ (.D(n1172),
	.CK(CLK),
	.Q(REGISTERS[65]));
   DFF_X1 REGISTERS_reg_29__0_ (.D(n1171),
	.CK(CLK),
	.Q(REGISTERS[64]));
   DFF_X1 REGISTERS_reg_30__31_ (.D(n1170),
	.CK(CLK),
	.Q(REGISTERS[63]));
   DFF_X1 REGISTERS_reg_30__30_ (.D(n1169),
	.CK(CLK),
	.Q(REGISTERS[62]));
   DFF_X1 REGISTERS_reg_30__29_ (.D(n1168),
	.CK(CLK),
	.Q(REGISTERS[61]));
   DFF_X1 REGISTERS_reg_30__28_ (.D(n1167),
	.CK(CLK),
	.Q(REGISTERS[60]));
   DFF_X1 REGISTERS_reg_30__27_ (.D(n1166),
	.CK(CLK),
	.Q(REGISTERS[59]));
   DFF_X1 REGISTERS_reg_30__26_ (.D(n1165),
	.CK(CLK),
	.Q(REGISTERS[58]));
   DFF_X1 REGISTERS_reg_30__25_ (.D(n1164),
	.CK(CLK),
	.Q(REGISTERS[57]));
   DFF_X1 REGISTERS_reg_30__24_ (.D(n1163),
	.CK(CLK),
	.Q(REGISTERS[56]));
   DFF_X1 REGISTERS_reg_30__23_ (.D(n1162),
	.CK(CLK),
	.Q(REGISTERS[55]));
   DFF_X1 REGISTERS_reg_30__22_ (.D(n1161),
	.CK(CLK),
	.Q(REGISTERS[54]));
   DFF_X1 REGISTERS_reg_30__21_ (.D(n1160),
	.CK(CLK),
	.Q(REGISTERS[53]));
   DFF_X1 REGISTERS_reg_30__20_ (.D(n1159),
	.CK(CLK),
	.Q(REGISTERS[52]));
   DFF_X1 REGISTERS_reg_30__19_ (.D(n1158),
	.CK(CLK),
	.Q(REGISTERS[51]));
   DFF_X1 REGISTERS_reg_30__18_ (.D(n1157),
	.CK(CLK),
	.Q(REGISTERS[50]));
   DFF_X1 REGISTERS_reg_30__17_ (.D(n1156),
	.CK(CLK),
	.Q(REGISTERS[49]));
   DFF_X1 REGISTERS_reg_30__16_ (.D(n1155),
	.CK(CLK),
	.Q(REGISTERS[48]));
   DFF_X1 REGISTERS_reg_30__15_ (.D(n1154),
	.CK(CLK),
	.Q(REGISTERS[47]));
   DFF_X1 REGISTERS_reg_30__14_ (.D(n1153),
	.CK(CLK),
	.Q(REGISTERS[46]));
   DFF_X1 REGISTERS_reg_30__13_ (.D(n1152),
	.CK(CLK),
	.Q(REGISTERS[45]));
   DFF_X1 REGISTERS_reg_30__12_ (.D(n1151),
	.CK(CLK),
	.Q(REGISTERS[44]));
   DFF_X1 REGISTERS_reg_30__11_ (.D(n1150),
	.CK(CLK),
	.Q(REGISTERS[43]));
   DFF_X1 REGISTERS_reg_30__10_ (.D(n1149),
	.CK(CLK),
	.Q(REGISTERS[42]));
   DFF_X1 REGISTERS_reg_30__9_ (.D(n1148),
	.CK(CLK),
	.Q(REGISTERS[41]));
   DFF_X1 REGISTERS_reg_30__8_ (.D(n1147),
	.CK(CLK),
	.Q(REGISTERS[40]));
   DFF_X1 REGISTERS_reg_30__7_ (.D(n1146),
	.CK(CLK),
	.Q(REGISTERS[39]));
   DFF_X1 REGISTERS_reg_30__6_ (.D(n1145),
	.CK(CLK),
	.Q(REGISTERS[38]));
   DFF_X1 REGISTERS_reg_30__5_ (.D(n1144),
	.CK(CLK),
	.Q(REGISTERS[37]));
   DFF_X1 REGISTERS_reg_30__4_ (.D(n1143),
	.CK(CLK),
	.Q(REGISTERS[36]));
   DFF_X1 REGISTERS_reg_30__3_ (.D(n1142),
	.CK(CLK),
	.Q(REGISTERS[35]));
   DFF_X1 REGISTERS_reg_30__2_ (.D(n1141),
	.CK(CLK),
	.Q(REGISTERS[34]));
   DFF_X1 REGISTERS_reg_30__1_ (.D(n1140),
	.CK(CLK),
	.Q(REGISTERS[33]));
   DFF_X1 REGISTERS_reg_30__0_ (.D(n1139),
	.CK(CLK),
	.Q(REGISTERS[32]));
   DFF_X1 REGISTERS_reg_31__31_ (.D(n1138),
	.CK(CLK),
	.Q(REGISTERS[31]));
   DFF_X1 REGISTERS_reg_31__30_ (.D(n1137),
	.CK(CLK),
	.Q(REGISTERS[30]));
   DFF_X1 REGISTERS_reg_31__29_ (.D(n1136),
	.CK(CLK),
	.Q(REGISTERS[29]));
   DFF_X1 REGISTERS_reg_31__28_ (.D(n1135),
	.CK(CLK),
	.Q(REGISTERS[28]));
   DFF_X1 REGISTERS_reg_31__27_ (.D(n1134),
	.CK(CLK),
	.Q(REGISTERS[27]));
   DFF_X1 REGISTERS_reg_31__26_ (.D(n1133),
	.CK(CLK),
	.Q(REGISTERS[26]));
   DFF_X1 REGISTERS_reg_31__25_ (.D(n1132),
	.CK(CLK),
	.Q(REGISTERS[25]));
   DFF_X1 REGISTERS_reg_31__24_ (.D(n1131),
	.CK(CLK),
	.Q(REGISTERS[24]));
   DFF_X1 REGISTERS_reg_31__23_ (.D(n1130),
	.CK(CLK),
	.Q(REGISTERS[23]));
   DFF_X1 REGISTERS_reg_31__22_ (.D(n1129),
	.CK(CLK),
	.Q(REGISTERS[22]));
   DFF_X1 REGISTERS_reg_31__21_ (.D(n1128),
	.CK(CLK),
	.Q(REGISTERS[21]));
   DFF_X1 REGISTERS_reg_31__20_ (.D(n1127),
	.CK(CLK),
	.Q(REGISTERS[20]));
   DFF_X1 REGISTERS_reg_31__19_ (.D(n1126),
	.CK(CLK),
	.Q(REGISTERS[19]));
   DFF_X1 REGISTERS_reg_31__18_ (.D(n1125),
	.CK(CLK),
	.Q(REGISTERS[18]));
   DFF_X1 REGISTERS_reg_31__17_ (.D(n1124),
	.CK(CLK),
	.Q(REGISTERS[17]));
   DFF_X1 REGISTERS_reg_31__16_ (.D(n1123),
	.CK(CLK),
	.Q(REGISTERS[16]));
   DFF_X1 REGISTERS_reg_31__15_ (.D(n1122),
	.CK(CLK),
	.Q(REGISTERS[15]));
   DFF_X1 REGISTERS_reg_31__14_ (.D(n1121),
	.CK(CLK),
	.Q(REGISTERS[14]));
   DFF_X1 REGISTERS_reg_31__13_ (.D(n1120),
	.CK(CLK),
	.Q(REGISTERS[13]));
   DFF_X1 REGISTERS_reg_31__12_ (.D(n1119),
	.CK(CLK),
	.Q(REGISTERS[12]));
   DFF_X1 REGISTERS_reg_31__11_ (.D(n1118),
	.CK(CLK),
	.Q(REGISTERS[11]));
   DFF_X1 REGISTERS_reg_31__10_ (.D(n1117),
	.CK(CLK),
	.Q(REGISTERS[10]));
   DFF_X1 REGISTERS_reg_31__9_ (.D(n1116),
	.CK(CLK),
	.Q(REGISTERS[9]));
   DFF_X1 REGISTERS_reg_31__8_ (.D(n1115),
	.CK(CLK),
	.Q(REGISTERS[8]));
   DFF_X1 REGISTERS_reg_31__7_ (.D(n1114),
	.CK(CLK),
	.Q(REGISTERS[7]));
   DFF_X1 REGISTERS_reg_31__6_ (.D(n1113),
	.CK(CLK),
	.Q(REGISTERS[6]));
   DFF_X1 REGISTERS_reg_31__5_ (.D(n1112),
	.CK(CLK),
	.Q(REGISTERS[5]));
   DFF_X1 REGISTERS_reg_31__4_ (.D(n1111),
	.CK(CLK),
	.Q(REGISTERS[4]));
   DFF_X1 REGISTERS_reg_31__3_ (.D(n1110),
	.CK(CLK),
	.Q(REGISTERS[3]));
   DFF_X1 REGISTERS_reg_31__2_ (.D(n1109),
	.CK(CLK),
	.Q(REGISTERS[2]));
   DFF_X1 REGISTERS_reg_31__1_ (.D(n1108),
	.CK(CLK),
	.Q(REGISTERS[1]));
   DFF_X1 REGISTERS_reg_31__0_ (.D(n1107),
	.CK(CLK),
	.Q(REGISTERS[0]));
   NAND3_X1 U2185 (.A1(ADD_WR[4]),
	.A2(ADD_WR[3]),
	.A3(WR),
	.ZN(n103));
   NAND3_X1 U2186 (.A1(ADD_WR[4]),
	.A2(n4037),
	.A3(WR),
	.ZN(n376));
   NAND3_X1 U2187 (.A1(ADD_WR[3]),
	.A2(n4020),
	.A3(WR),
	.ZN(n641));
   NAND3_X1 U2188 (.A1(n4039),
	.A2(n4038),
	.A3(n4040),
	.ZN(n342));
   NAND3_X1 U2189 (.A1(ADD_WR[1]),
	.A2(ADD_WR[0]),
	.A3(ADD_WR[2]),
	.ZN(n104));
   NAND3_X1 U2190 (.A1(ADD_WR[1]),
	.A2(n4040),
	.A3(ADD_WR[2]),
	.ZN(n138));
   NAND3_X1 U2191 (.A1(ADD_WR[0]),
	.A2(n4039),
	.A3(ADD_WR[2]),
	.ZN(n172));
   NAND3_X1 U2192 (.A1(n4040),
	.A2(n4039),
	.A3(ADD_WR[2]),
	.ZN(n206));
   NAND3_X1 U2193 (.A1(ADD_WR[0]),
	.A2(n4038),
	.A3(ADD_WR[1]),
	.ZN(n240));
   NAND3_X1 U2194 (.A1(n4040),
	.A2(n4038),
	.A3(ADD_WR[1]),
	.ZN(n274));
   NAND3_X1 U2195 (.A1(n4037),
	.A2(n4020),
	.A3(WR),
	.ZN(n906));
   NAND3_X1 U2196 (.A1(n4039),
	.A2(n4038),
	.A3(ADD_WR[0]),
	.ZN(n308));
   AND2_X1 U436 (.A1(N55),
	.A2(n1106),
	.ZN(OUT1[7]));
   AND2_X1 U437 (.A1(N56),
	.A2(n1106),
	.ZN(OUT1[6]));
   AND2_X1 U438 (.A1(N57),
	.A2(n1106),
	.ZN(OUT1[5]));
   AND2_X1 U439 (.A1(N58),
	.A2(n1106),
	.ZN(OUT1[4]));
   AND2_X1 U440 (.A1(N59),
	.A2(n1106),
	.ZN(OUT1[3]));
   AND2_X1 U441 (.A1(N60),
	.A2(n1106),
	.ZN(OUT1[2]));
   AND2_X1 U442 (.A1(N61),
	.A2(n1106),
	.ZN(OUT1[1]));
   AND2_X1 U443 (.A1(N62),
	.A2(n1106),
	.ZN(OUT1[0]));
   AND2_X1 U444 (.A1(N39),
	.A2(n1106),
	.ZN(OUT1[23]));
   AND2_X1 U445 (.A1(N40),
	.A2(n1106),
	.ZN(OUT1[22]));
   AND2_X1 U446 (.A1(N41),
	.A2(n1106),
	.ZN(OUT1[21]));
   AND2_X1 U447 (.A1(N42),
	.A2(n1106),
	.ZN(OUT1[20]));
   AND2_X1 U448 (.A1(N31),
	.A2(n1106),
	.ZN(OUT1[31]));
   AND2_X1 U449 (.A1(N32),
	.A2(n1106),
	.ZN(OUT1[30]));
   AND2_X1 U450 (.A1(N33),
	.A2(n1106),
	.ZN(OUT1[29]));
   AND2_X1 U451 (.A1(N34),
	.A2(n1106),
	.ZN(OUT1[28]));
   AND2_X1 U452 (.A1(N35),
	.A2(n1106),
	.ZN(OUT1[27]));
   AND2_X1 U453 (.A1(N36),
	.A2(n1106),
	.ZN(OUT1[26]));
   AND2_X1 U454 (.A1(N37),
	.A2(n1106),
	.ZN(OUT1[25]));
   AND2_X1 U455 (.A1(N38),
	.A2(n1106),
	.ZN(OUT1[24]));
   AND2_X1 U456 (.A1(N43),
	.A2(n1106),
	.ZN(OUT1[19]));
   AND2_X1 U457 (.A1(N44),
	.A2(n1106),
	.ZN(OUT1[18]));
   AND2_X1 U458 (.A1(N45),
	.A2(n1106),
	.ZN(OUT1[17]));
   AND2_X1 U459 (.A1(N46),
	.A2(n1106),
	.ZN(OUT1[16]));
   AND2_X1 U460 (.A1(N47),
	.A2(n1106),
	.ZN(OUT1[15]));
   AND2_X1 U461 (.A1(N48),
	.A2(n1106),
	.ZN(OUT1[14]));
   AND2_X1 U462 (.A1(N49),
	.A2(n1106),
	.ZN(OUT1[13]));
   AND2_X1 U463 (.A1(N50),
	.A2(n1106),
	.ZN(OUT1[12]));
   AND2_X1 U464 (.A1(N51),
	.A2(n1106),
	.ZN(OUT1[11]));
   AND2_X1 U465 (.A1(N52),
	.A2(n1106),
	.ZN(OUT1[10]));
   AND2_X1 U466 (.A1(N53),
	.A2(n1106),
	.ZN(OUT1[9]));
   AND2_X1 U467 (.A1(N54),
	.A2(n1106),
	.ZN(OUT1[8]));
   AND2_X1 U468 (.A1(N104),
	.A2(n1105),
	.ZN(OUT2[23]));
   AND2_X1 U469 (.A1(N105),
	.A2(n1105),
	.ZN(OUT2[22]));
   AND2_X1 U470 (.A1(N106),
	.A2(n1105),
	.ZN(OUT2[21]));
   AND2_X1 U471 (.A1(N107),
	.A2(n1105),
	.ZN(OUT2[20]));
   AND2_X1 U472 (.A1(N96),
	.A2(n1105),
	.ZN(OUT2[31]));
   AND2_X1 U473 (.A1(N97),
	.A2(n1105),
	.ZN(OUT2[30]));
   AND2_X1 U474 (.A1(N98),
	.A2(n1105),
	.ZN(OUT2[29]));
   AND2_X1 U475 (.A1(N99),
	.A2(n1105),
	.ZN(OUT2[28]));
   AND2_X1 U476 (.A1(N100),
	.A2(n1105),
	.ZN(OUT2[27]));
   AND2_X1 U477 (.A1(N101),
	.A2(n1105),
	.ZN(OUT2[26]));
   AND2_X1 U478 (.A1(N102),
	.A2(n1105),
	.ZN(OUT2[25]));
   AND2_X1 U479 (.A1(N103),
	.A2(n1105),
	.ZN(OUT2[24]));
   AND2_X1 U480 (.A1(N108),
	.A2(n1105),
	.ZN(OUT2[19]));
   AND2_X1 U481 (.A1(N109),
	.A2(n1105),
	.ZN(OUT2[18]));
   AND2_X1 U482 (.A1(N110),
	.A2(n1105),
	.ZN(OUT2[17]));
   AND2_X1 U483 (.A1(N111),
	.A2(n1105),
	.ZN(OUT2[16]));
   AND2_X1 U484 (.A1(N112),
	.A2(n1105),
	.ZN(OUT2[15]));
   AND2_X1 U485 (.A1(N113),
	.A2(n1105),
	.ZN(OUT2[14]));
   AND2_X1 U486 (.A1(N114),
	.A2(n1105),
	.ZN(OUT2[13]));
   AND2_X1 U487 (.A1(N115),
	.A2(n1105),
	.ZN(OUT2[12]));
   AND2_X1 U488 (.A1(N116),
	.A2(n1105),
	.ZN(OUT2[11]));
   AND2_X1 U489 (.A1(N117),
	.A2(n1105),
	.ZN(OUT2[10]));
   AND2_X1 U490 (.A1(N118),
	.A2(n1105),
	.ZN(OUT2[9]));
   AND2_X1 U491 (.A1(N119),
	.A2(n1105),
	.ZN(OUT2[8]));
   AND2_X1 U492 (.A1(N120),
	.A2(n1105),
	.ZN(OUT2[7]));
   AND2_X1 U493 (.A1(N121),
	.A2(n1105),
	.ZN(OUT2[6]));
   AND2_X1 U494 (.A1(N122),
	.A2(n1105),
	.ZN(OUT2[5]));
   AND2_X1 U495 (.A1(N123),
	.A2(n1105),
	.ZN(OUT2[4]));
   AND2_X1 U496 (.A1(N124),
	.A2(n1105),
	.ZN(OUT2[3]));
   AND2_X1 U497 (.A1(N125),
	.A2(n1105),
	.ZN(OUT2[2]));
   AND2_X1 U498 (.A1(N126),
	.A2(n1105),
	.ZN(OUT2[1]));
   AND2_X1 U499 (.A1(N127),
	.A2(n1105),
	.ZN(OUT2[0]));
   AND2_X2 U540 (.A1(RD1),
	.A2(ENABLE),
	.ZN(n1106));
   AND2_X2 U541 (.A1(RD2),
	.A2(ENABLE),
	.ZN(n1105));
   NAND2_X2 U549 (.A1(DATAIN[0]),
	.A2(n4041),
	.ZN(n38));
   NAND2_X2 U550 (.A1(DATAIN[1]),
	.A2(n4041),
	.ZN(n40));
   NAND2_X2 U551 (.A1(DATAIN[2]),
	.A2(n4041),
	.ZN(n42));
   NAND2_X2 U552 (.A1(DATAIN[3]),
	.A2(n4041),
	.ZN(n44));
   NAND2_X2 U553 (.A1(DATAIN[4]),
	.A2(n4041),
	.ZN(n46));
   NAND2_X2 U554 (.A1(DATAIN[6]),
	.A2(n4041),
	.ZN(n50));
   NAND2_X2 U555 (.A1(DATAIN[8]),
	.A2(n4041),
	.ZN(n54));
   NAND2_X2 U556 (.A1(DATAIN[9]),
	.A2(n4041),
	.ZN(n56));
   NAND2_X2 U557 (.A1(DATAIN[10]),
	.A2(n4041),
	.ZN(n58));
   NAND2_X2 U558 (.A1(DATAIN[12]),
	.A2(n4041),
	.ZN(n62));
   NAND2_X2 U559 (.A1(DATAIN[14]),
	.A2(n4041),
	.ZN(n66));
   NAND2_X2 U560 (.A1(DATAIN[16]),
	.A2(n4041),
	.ZN(n70));
   NAND2_X2 U561 (.A1(DATAIN[18]),
	.A2(n4041),
	.ZN(n74));
   NAND2_X2 U562 (.A1(DATAIN[19]),
	.A2(n4041),
	.ZN(n76));
   NAND2_X2 U563 (.A1(DATAIN[20]),
	.A2(n4041),
	.ZN(n78));
   NAND2_X2 U564 (.A1(DATAIN[22]),
	.A2(n4041),
	.ZN(n82));
   NAND2_X2 U565 (.A1(DATAIN[24]),
	.A2(n4041),
	.ZN(n86));
   NAND2_X2 U566 (.A1(DATAIN[25]),
	.A2(n4041),
	.ZN(n88));
   NAND2_X2 U567 (.A1(DATAIN[26]),
	.A2(n4041),
	.ZN(n90));
   NAND2_X2 U568 (.A1(DATAIN[27]),
	.A2(n4041),
	.ZN(n92));
   NAND2_X2 U569 (.A1(DATAIN[28]),
	.A2(n4041),
	.ZN(n94));
   NAND2_X2 U570 (.A1(DATAIN[29]),
	.A2(n4041),
	.ZN(n96));
   NAND2_X2 U571 (.A1(DATAIN[30]),
	.A2(n4041),
	.ZN(n98));
   NAND2_X2 U572 (.A1(DATAIN[31]),
	.A2(n4041),
	.ZN(n100));
   INV_X2 U573 (.A(n375),
	.ZN(n4036));
   OAI21_X1 U574 (.A(n4041),
	.B1(n104),
	.B2(n376),
	.ZN(n375));
   INV_X2 U575 (.A(n409),
	.ZN(n4035));
   OAI21_X1 U576 (.A(FE_OFN18_n4041),
	.B1(n138),
	.B2(n376),
	.ZN(n409));
   INV_X1 U577 (.A(n442),
	.ZN(n4034));
   OAI21_X1 U578 (.A(FE_OFN18_n4041),
	.B1(n172),
	.B2(n376),
	.ZN(n442));
   INV_X1 U579 (.A(n475),
	.ZN(n4033));
   OAI21_X1 U580 (.A(FE_OFN18_n4041),
	.B1(n206),
	.B2(n376),
	.ZN(n475));
   INV_X2 U581 (.A(n508),
	.ZN(n4032));
   OAI21_X1 U582 (.A(n4041),
	.B1(n240),
	.B2(n376),
	.ZN(n508));
   INV_X1 U583 (.A(n541),
	.ZN(n4031));
   OAI21_X1 U584 (.A(n4041),
	.B1(n274),
	.B2(n376),
	.ZN(n541));
   INV_X2 U585 (.A(n574),
	.ZN(n4030));
   OAI21_X1 U586 (.A(n4041),
	.B1(n308),
	.B2(n376),
	.ZN(n574));
   INV_X2 U587 (.A(n607),
	.ZN(n4029));
   OAI21_X1 U588 (.A(n4041),
	.B1(n342),
	.B2(n376),
	.ZN(n607));
   INV_X2 U589 (.A(n640),
	.ZN(n4019));
   OAI21_X1 U590 (.A(FE_OFN18_n4041),
	.B1(n104),
	.B2(n641),
	.ZN(n640));
   INV_X1 U591 (.A(n674),
	.ZN(n4018));
   OAI21_X1 U592 (.A(FE_OFN18_n4041),
	.B1(n138),
	.B2(n641),
	.ZN(n674));
   INV_X2 U593 (.A(n707),
	.ZN(n4017));
   OAI21_X1 U594 (.A(FE_OFN18_n4041),
	.B1(n172),
	.B2(n641),
	.ZN(n707));
   INV_X1 U595 (.A(n740),
	.ZN(n4016));
   OAI21_X1 U596 (.A(FE_OFN18_n4041),
	.B1(n206),
	.B2(n641),
	.ZN(n740));
   INV_X2 U597 (.A(n773),
	.ZN(n4015));
   OAI21_X1 U598 (.A(FE_OFN18_n4041),
	.B1(n240),
	.B2(n641),
	.ZN(n773));
   INV_X2 U599 (.A(n806),
	.ZN(n4014));
   OAI21_X1 U600 (.A(FE_OFN18_n4041),
	.B1(n274),
	.B2(n641),
	.ZN(n806));
   INV_X2 U601 (.A(n839),
	.ZN(n4013));
   OAI21_X1 U602 (.A(FE_OFN18_n4041),
	.B1(n308),
	.B2(n641),
	.ZN(n839));
   INV_X2 U603 (.A(n872),
	.ZN(n4012));
   OAI21_X1 U604 (.A(FE_OFN18_n4041),
	.B1(n342),
	.B2(n641),
	.ZN(n872));
   NAND2_X2 U605 (.A1(DATAIN[5]),
	.A2(n4041),
	.ZN(n48));
   NAND2_X2 U606 (.A1(DATAIN[7]),
	.A2(n4041),
	.ZN(n52));
   NAND2_X2 U607 (.A1(DATAIN[11]),
	.A2(n4041),
	.ZN(n60));
   NAND2_X2 U608 (.A1(DATAIN[13]),
	.A2(n4041),
	.ZN(n64));
   NAND2_X2 U609 (.A1(DATAIN[15]),
	.A2(n4041),
	.ZN(n68));
   NAND2_X2 U610 (.A1(DATAIN[17]),
	.A2(n4041),
	.ZN(n72));
   NAND2_X2 U611 (.A1(DATAIN[21]),
	.A2(n4041),
	.ZN(n80));
   NAND2_X2 U612 (.A1(DATAIN[23]),
	.A2(n4041),
	.ZN(n84));
   INV_X2 U613 (.A(n905),
	.ZN(n4011));
   OAI21_X1 U614 (.A(FE_OFN18_n4041),
	.B1(n104),
	.B2(n906),
	.ZN(n905));
   INV_X2 U615 (.A(n939),
	.ZN(n4010));
   OAI21_X1 U616 (.A(FE_OFN18_n4041),
	.B1(n138),
	.B2(n906),
	.ZN(n939));
   INV_X2 U617 (.A(n972),
	.ZN(n4009));
   OAI21_X1 U618 (.A(FE_OFN18_n4041),
	.B1(n172),
	.B2(n906),
	.ZN(n972));
   INV_X2 U619 (.A(n1005),
	.ZN(n4008));
   OAI21_X1 U620 (.A(FE_OFN18_n4041),
	.B1(n206),
	.B2(n906),
	.ZN(n1005));
   INV_X2 U621 (.A(n1038),
	.ZN(n4007));
   OAI21_X1 U622 (.A(FE_OFN18_n4041),
	.B1(n240),
	.B2(n906),
	.ZN(n1038));
   INV_X1 U623 (.A(n1071),
	.ZN(n4006));
   OAI21_X1 U624 (.A(FE_OFN18_n4041),
	.B1(n274),
	.B2(n906),
	.ZN(n1071));
   INV_X2 U625 (.A(n1104),
	.ZN(n4005));
   OAI21_X1 U626 (.A(FE_OFN18_n4041),
	.B1(n308),
	.B2(n906),
	.ZN(n1104));
   INV_X2 U627 (.A(n102),
	.ZN(n4028));
   OAI21_X1 U628 (.A(n4041),
	.B1(n103),
	.B2(n104),
	.ZN(n102));
   INV_X2 U629 (.A(n137),
	.ZN(n4027));
   OAI21_X1 U630 (.A(n4041),
	.B1(n103),
	.B2(n138),
	.ZN(n137));
   INV_X2 U631 (.A(n171),
	.ZN(n4026));
   OAI21_X1 U632 (.A(FE_OFN18_n4041),
	.B1(n103),
	.B2(n172),
	.ZN(n171));
   INV_X1 U633 (.A(n205),
	.ZN(n4025));
   OAI21_X1 U634 (.A(FE_OFN18_n4041),
	.B1(n103),
	.B2(n206),
	.ZN(n205));
   INV_X2 U635 (.A(n239),
	.ZN(n4024));
   OAI21_X1 U636 (.A(n4041),
	.B1(n103),
	.B2(n240),
	.ZN(n239));
   INV_X2 U637 (.A(n273),
	.ZN(n4023));
   OAI21_X1 U638 (.A(FE_OFN18_n4041),
	.B1(n103),
	.B2(n274),
	.ZN(n273));
   INV_X2 U639 (.A(n307),
	.ZN(n4022));
   OAI21_X1 U640 (.A(FE_OFN18_n4041),
	.B1(n103),
	.B2(n308),
	.ZN(n307));
   INV_X2 U641 (.A(n341),
	.ZN(n4021));
   OAI21_X1 U642 (.A(n4041),
	.B1(n103),
	.B2(n342),
	.ZN(n341));
   INV_X1 U643 (.A(ADD_RD1[0]),
	.ZN(n2782));
   INV_X1 U644 (.A(ADD_RD2[0]),
	.ZN(n3590));
   INV_X1 U645 (.A(ADD_RD1[2]),
	.ZN(n2784));
   INV_X1 U646 (.A(ADD_RD2[2]),
	.ZN(n3592));
   INV_X1 U647 (.A(ADD_RD1[1]),
	.ZN(n2783));
   INV_X1 U648 (.A(ADD_RD2[1]),
	.ZN(n3591));
   INV_X1 U649 (.A(ADD_RD1[3]),
	.ZN(n2785));
   INV_X1 U650 (.A(ADD_RD2[3]),
	.ZN(n3593));
   INV_X1 U651 (.A(ADD_WR[2]),
	.ZN(n4038));
   OAI21_X1 U652 (.A(n53),
	.B1(FE_OFN75_n4028),
	.B2(n52),
	.ZN(n1114));
   NAND2_X1 U653 (.A1(REGISTERS[7]),
	.A2(FE_OFN75_n4028),
	.ZN(n53));
   OAI21_X1 U654 (.A(n55),
	.B1(n4028),
	.B2(n54),
	.ZN(n1115));
   NAND2_X1 U655 (.A1(REGISTERS[8]),
	.A2(n4028),
	.ZN(n55));
   OAI21_X1 U656 (.A(n57),
	.B1(FE_OFN75_n4028),
	.B2(n56),
	.ZN(n1116));
   NAND2_X1 U657 (.A1(REGISTERS[9]),
	.A2(FE_OFN75_n4028),
	.ZN(n57));
   OAI21_X1 U658 (.A(n59),
	.B1(n4028),
	.B2(n58),
	.ZN(n1117));
   NAND2_X1 U659 (.A1(REGISTERS[10]),
	.A2(n4028),
	.ZN(n59));
   OAI21_X1 U660 (.A(n61),
	.B1(FE_OFN75_n4028),
	.B2(n60),
	.ZN(n1118));
   NAND2_X1 U661 (.A1(REGISTERS[11]),
	.A2(FE_OFN75_n4028),
	.ZN(n61));
   OAI21_X1 U662 (.A(n63),
	.B1(n4028),
	.B2(n62),
	.ZN(n1119));
   NAND2_X1 U663 (.A1(REGISTERS[12]),
	.A2(n4028),
	.ZN(n63));
   OAI21_X1 U664 (.A(n67),
	.B1(FE_OFN75_n4028),
	.B2(n66),
	.ZN(n1121));
   NAND2_X1 U665 (.A1(REGISTERS[14]),
	.A2(FE_OFN75_n4028),
	.ZN(n67));
   OAI21_X1 U666 (.A(n69),
	.B1(n4028),
	.B2(n68),
	.ZN(n1122));
   NAND2_X1 U667 (.A1(REGISTERS[15]),
	.A2(n4028),
	.ZN(n69));
   OAI21_X1 U668 (.A(n112),
	.B1(FE_OFN89_n4027),
	.B2(n52),
	.ZN(n1146));
   NAND2_X1 U669 (.A1(REGISTERS[39]),
	.A2(FE_OFN89_n4027),
	.ZN(n112));
   OAI21_X1 U670 (.A(n113),
	.B1(n4027),
	.B2(n54),
	.ZN(n1147));
   NAND2_X1 U671 (.A1(REGISTERS[40]),
	.A2(n4027),
	.ZN(n113));
   OAI21_X1 U672 (.A(n114),
	.B1(FE_OFN89_n4027),
	.B2(n56),
	.ZN(n1148));
   NAND2_X1 U673 (.A1(REGISTERS[41]),
	.A2(FE_OFN89_n4027),
	.ZN(n114));
   OAI21_X1 U674 (.A(n115),
	.B1(n4027),
	.B2(n58),
	.ZN(n1149));
   NAND2_X1 U675 (.A1(REGISTERS[42]),
	.A2(n4027),
	.ZN(n115));
   OAI21_X1 U676 (.A(n116),
	.B1(FE_OFN89_n4027),
	.B2(n60),
	.ZN(n1150));
   NAND2_X1 U677 (.A1(REGISTERS[43]),
	.A2(FE_OFN89_n4027),
	.ZN(n116));
   OAI21_X1 U678 (.A(n117),
	.B1(n4027),
	.B2(n62),
	.ZN(n1151));
   NAND2_X1 U679 (.A1(REGISTERS[44]),
	.A2(n4027),
	.ZN(n117));
   OAI21_X1 U680 (.A(n119),
	.B1(FE_OFN89_n4027),
	.B2(n66),
	.ZN(n1153));
   NAND2_X1 U681 (.A1(REGISTERS[46]),
	.A2(FE_OFN89_n4027),
	.ZN(n119));
   OAI21_X1 U682 (.A(n120),
	.B1(FE_OFN89_n4027),
	.B2(n68),
	.ZN(n1154));
   NAND2_X1 U683 (.A1(REGISTERS[47]),
	.A2(n4027),
	.ZN(n120));
   OAI21_X1 U684 (.A(n146),
	.B1(FE_OFN77_n4026),
	.B2(n52),
	.ZN(n1178));
   NAND2_X1 U685 (.A1(REGISTERS[71]),
	.A2(FE_OFN77_n4026),
	.ZN(n146));
   OAI21_X1 U686 (.A(n147),
	.B1(n4026),
	.B2(n54),
	.ZN(n1179));
   NAND2_X1 U687 (.A1(REGISTERS[72]),
	.A2(n4026),
	.ZN(n147));
   OAI21_X1 U688 (.A(n148),
	.B1(FE_OFN77_n4026),
	.B2(n56),
	.ZN(n1180));
   NAND2_X1 U689 (.A1(REGISTERS[73]),
	.A2(FE_OFN77_n4026),
	.ZN(n148));
   OAI21_X1 U690 (.A(n149),
	.B1(n4026),
	.B2(n58),
	.ZN(n1181));
   NAND2_X1 U691 (.A1(REGISTERS[74]),
	.A2(n4026),
	.ZN(n149));
   OAI21_X1 U692 (.A(n150),
	.B1(FE_OFN77_n4026),
	.B2(n60),
	.ZN(n1182));
   NAND2_X1 U693 (.A1(REGISTERS[75]),
	.A2(FE_OFN77_n4026),
	.ZN(n150));
   OAI21_X1 U694 (.A(n151),
	.B1(n4026),
	.B2(n62),
	.ZN(n1183));
   NAND2_X1 U695 (.A1(REGISTERS[76]),
	.A2(n4026),
	.ZN(n151));
   OAI21_X1 U696 (.A(n153),
	.B1(FE_OFN77_n4026),
	.B2(n66),
	.ZN(n1185));
   NAND2_X1 U697 (.A1(REGISTERS[78]),
	.A2(FE_OFN77_n4026),
	.ZN(n153));
   OAI21_X1 U698 (.A(n154),
	.B1(n4026),
	.B2(n68),
	.ZN(n1186));
   NAND2_X1 U699 (.A1(REGISTERS[79]),
	.A2(n4026),
	.ZN(n154));
   OAI21_X1 U700 (.A(n180),
	.B1(FE_OFN69_n4025),
	.B2(n52),
	.ZN(n1210));
   NAND2_X1 U701 (.A1(REGISTERS[103]),
	.A2(FE_OFN69_n4025),
	.ZN(n180));
   OAI21_X1 U702 (.A(n181),
	.B1(FE_OFN69_n4025),
	.B2(n54),
	.ZN(n1211));
   NAND2_X1 U703 (.A1(REGISTERS[104]),
	.A2(FE_OFN69_n4025),
	.ZN(n181));
   OAI21_X1 U704 (.A(n182),
	.B1(n4025),
	.B2(n56),
	.ZN(n1212));
   NAND2_X1 U705 (.A1(REGISTERS[105]),
	.A2(n4025),
	.ZN(n182));
   OAI21_X1 U706 (.A(n183),
	.B1(n4025),
	.B2(n58),
	.ZN(n1213));
   NAND2_X1 U707 (.A1(REGISTERS[106]),
	.A2(n4025),
	.ZN(n183));
   OAI21_X1 U708 (.A(n184),
	.B1(FE_OFN69_n4025),
	.B2(n60),
	.ZN(n1214));
   NAND2_X1 U709 (.A1(REGISTERS[107]),
	.A2(FE_OFN69_n4025),
	.ZN(n184));
   OAI21_X1 U710 (.A(n185),
	.B1(n4025),
	.B2(n62),
	.ZN(n1215));
   NAND2_X1 U711 (.A1(REGISTERS[108]),
	.A2(n4025),
	.ZN(n185));
   OAI21_X1 U712 (.A(n187),
	.B1(FE_OFN69_n4025),
	.B2(n66),
	.ZN(n1217));
   NAND2_X1 U713 (.A1(REGISTERS[110]),
	.A2(FE_OFN69_n4025),
	.ZN(n187));
   OAI21_X1 U714 (.A(n188),
	.B1(n4025),
	.B2(n68),
	.ZN(n1218));
   NAND2_X1 U715 (.A1(REGISTERS[111]),
	.A2(n4025),
	.ZN(n188));
   OAI21_X1 U716 (.A(n207),
	.B1(FE_OFN83_n4024),
	.B2(n38),
	.ZN(n1235));
   NAND2_X1 U717 (.A1(REGISTERS[128]),
	.A2(FE_OFN83_n4024),
	.ZN(n207));
   OAI21_X1 U718 (.A(n209),
	.B1(FE_OFN83_n4024),
	.B2(n42),
	.ZN(n1237));
   NAND2_X1 U719 (.A1(REGISTERS[130]),
	.A2(FE_OFN83_n4024),
	.ZN(n209));
   OAI21_X1 U720 (.A(n212),
	.B1(FE_OFN83_n4024),
	.B2(n48),
	.ZN(n1240));
   NAND2_X1 U721 (.A1(REGISTERS[133]),
	.A2(FE_OFN83_n4024),
	.ZN(n212));
   OAI21_X1 U722 (.A(n213),
	.B1(n4024),
	.B2(n50),
	.ZN(n1241));
   NAND2_X1 U723 (.A1(REGISTERS[134]),
	.A2(n4024),
	.ZN(n213));
   OAI21_X1 U724 (.A(n214),
	.B1(FE_OFN83_n4024),
	.B2(n52),
	.ZN(n1242));
   NAND2_X1 U725 (.A1(REGISTERS[135]),
	.A2(FE_OFN83_n4024),
	.ZN(n214));
   OAI21_X1 U726 (.A(n215),
	.B1(n4024),
	.B2(n54),
	.ZN(n1243));
   NAND2_X1 U727 (.A1(REGISTERS[136]),
	.A2(n4024),
	.ZN(n215));
   OAI21_X1 U728 (.A(n216),
	.B1(FE_OFN83_n4024),
	.B2(n56),
	.ZN(n1244));
   NAND2_X1 U729 (.A1(REGISTERS[137]),
	.A2(FE_OFN83_n4024),
	.ZN(n216));
   OAI21_X1 U730 (.A(n217),
	.B1(n4024),
	.B2(n58),
	.ZN(n1245));
   NAND2_X1 U731 (.A1(REGISTERS[138]),
	.A2(n4024),
	.ZN(n217));
   OAI21_X1 U732 (.A(n218),
	.B1(FE_OFN83_n4024),
	.B2(n60),
	.ZN(n1246));
   NAND2_X1 U733 (.A1(REGISTERS[139]),
	.A2(FE_OFN83_n4024),
	.ZN(n218));
   OAI21_X1 U734 (.A(n219),
	.B1(n4024),
	.B2(n62),
	.ZN(n1247));
   NAND2_X1 U735 (.A1(REGISTERS[140]),
	.A2(n4024),
	.ZN(n219));
   OAI21_X1 U736 (.A(n220),
	.B1(n4024),
	.B2(n64),
	.ZN(n1248));
   NAND2_X1 U737 (.A1(REGISTERS[141]),
	.A2(n4024),
	.ZN(n220));
   OAI21_X1 U738 (.A(n221),
	.B1(FE_OFN83_n4024),
	.B2(n66),
	.ZN(n1249));
   NAND2_X1 U739 (.A1(REGISTERS[142]),
	.A2(FE_OFN83_n4024),
	.ZN(n221));
   OAI21_X1 U740 (.A(n222),
	.B1(n4024),
	.B2(n68),
	.ZN(n1250));
   NAND2_X1 U741 (.A1(REGISTERS[143]),
	.A2(n4024),
	.ZN(n222));
   OAI21_X1 U742 (.A(n223),
	.B1(FE_OFN83_n4024),
	.B2(n70),
	.ZN(n1251));
   NAND2_X1 U743 (.A1(REGISTERS[144]),
	.A2(FE_OFN83_n4024),
	.ZN(n223));
   OAI21_X1 U744 (.A(n224),
	.B1(FE_OFN83_n4024),
	.B2(n72),
	.ZN(n1252));
   NAND2_X1 U745 (.A1(REGISTERS[145]),
	.A2(FE_OFN83_n4024),
	.ZN(n224));
   OAI21_X1 U746 (.A(n225),
	.B1(n4024),
	.B2(n74),
	.ZN(n1253));
   NAND2_X1 U747 (.A1(REGISTERS[146]),
	.A2(n4024),
	.ZN(n225));
   OAI21_X1 U748 (.A(n226),
	.B1(FE_OFN83_n4024),
	.B2(n76),
	.ZN(n1254));
   NAND2_X1 U749 (.A1(REGISTERS[147]),
	.A2(FE_OFN83_n4024),
	.ZN(n226));
   OAI21_X1 U750 (.A(n227),
	.B1(n4024),
	.B2(n78),
	.ZN(n1255));
   NAND2_X1 U751 (.A1(REGISTERS[148]),
	.A2(n4024),
	.ZN(n227));
   OAI21_X1 U752 (.A(n228),
	.B1(FE_OFN83_n4024),
	.B2(n80),
	.ZN(n1256));
   NAND2_X1 U753 (.A1(REGISTERS[149]),
	.A2(FE_OFN83_n4024),
	.ZN(n228));
   OAI21_X1 U754 (.A(n229),
	.B1(FE_OFN83_n4024),
	.B2(n82),
	.ZN(n1257));
   NAND2_X1 U755 (.A1(REGISTERS[150]),
	.A2(FE_OFN83_n4024),
	.ZN(n229));
   OAI21_X1 U756 (.A(n230),
	.B1(FE_OFN83_n4024),
	.B2(n84),
	.ZN(n1258));
   NAND2_X1 U757 (.A1(REGISTERS[151]),
	.A2(FE_OFN83_n4024),
	.ZN(n230));
   OAI21_X1 U758 (.A(n231),
	.B1(n4024),
	.B2(n86),
	.ZN(n1259));
   NAND2_X1 U759 (.A1(REGISTERS[152]),
	.A2(n4024),
	.ZN(n231));
   OAI21_X1 U760 (.A(n232),
	.B1(FE_OFN83_n4024),
	.B2(n88),
	.ZN(n1260));
   NAND2_X1 U761 (.A1(REGISTERS[153]),
	.A2(FE_OFN83_n4024),
	.ZN(n232));
   OAI21_X1 U762 (.A(n233),
	.B1(n4024),
	.B2(n90),
	.ZN(n1261));
   NAND2_X1 U763 (.A1(REGISTERS[154]),
	.A2(n4024),
	.ZN(n233));
   OAI21_X1 U764 (.A(n234),
	.B1(FE_OFN83_n4024),
	.B2(n92),
	.ZN(n1262));
   NAND2_X1 U765 (.A1(REGISTERS[155]),
	.A2(FE_OFN83_n4024),
	.ZN(n234));
   OAI21_X1 U766 (.A(n235),
	.B1(FE_OFN83_n4024),
	.B2(n94),
	.ZN(n1263));
   NAND2_X1 U767 (.A1(REGISTERS[156]),
	.A2(FE_OFN83_n4024),
	.ZN(n235));
   OAI21_X1 U768 (.A(n248),
	.B1(FE_OFN79_n4023),
	.B2(n52),
	.ZN(n1274));
   NAND2_X1 U769 (.A1(REGISTERS[167]),
	.A2(FE_OFN79_n4023),
	.ZN(n248));
   OAI21_X1 U770 (.A(n249),
	.B1(n4023),
	.B2(n54),
	.ZN(n1275));
   NAND2_X1 U771 (.A1(REGISTERS[168]),
	.A2(n4023),
	.ZN(n249));
   OAI21_X1 U772 (.A(n250),
	.B1(FE_OFN79_n4023),
	.B2(n56),
	.ZN(n1276));
   NAND2_X1 U773 (.A1(REGISTERS[169]),
	.A2(FE_OFN79_n4023),
	.ZN(n250));
   OAI21_X1 U774 (.A(n251),
	.B1(n4023),
	.B2(n58),
	.ZN(n1277));
   NAND2_X1 U775 (.A1(REGISTERS[170]),
	.A2(n4023),
	.ZN(n251));
   OAI21_X1 U776 (.A(n252),
	.B1(FE_OFN79_n4023),
	.B2(n60),
	.ZN(n1278));
   NAND2_X1 U777 (.A1(REGISTERS[171]),
	.A2(FE_OFN79_n4023),
	.ZN(n252));
   OAI21_X1 U778 (.A(n253),
	.B1(n4023),
	.B2(n62),
	.ZN(n1279));
   NAND2_X1 U779 (.A1(REGISTERS[172]),
	.A2(n4023),
	.ZN(n253));
   OAI21_X1 U780 (.A(n255),
	.B1(FE_OFN79_n4023),
	.B2(n66),
	.ZN(n1281));
   NAND2_X1 U781 (.A1(REGISTERS[174]),
	.A2(FE_OFN79_n4023),
	.ZN(n255));
   OAI21_X1 U782 (.A(n256),
	.B1(n4023),
	.B2(n68),
	.ZN(n1282));
   NAND2_X1 U783 (.A1(REGISTERS[175]),
	.A2(n4023),
	.ZN(n256));
   OAI21_X1 U784 (.A(n282),
	.B1(FE_OFN85_n4022),
	.B2(n52),
	.ZN(n1306));
   NAND2_X1 U785 (.A1(REGISTERS[199]),
	.A2(FE_OFN85_n4022),
	.ZN(n282));
   OAI21_X1 U786 (.A(n283),
	.B1(n4022),
	.B2(n54),
	.ZN(n1307));
   NAND2_X1 U787 (.A1(REGISTERS[200]),
	.A2(n4022),
	.ZN(n283));
   OAI21_X1 U788 (.A(n284),
	.B1(FE_OFN85_n4022),
	.B2(n56),
	.ZN(n1308));
   NAND2_X1 U789 (.A1(REGISTERS[201]),
	.A2(FE_OFN85_n4022),
	.ZN(n284));
   OAI21_X1 U790 (.A(n285),
	.B1(n4022),
	.B2(n58),
	.ZN(n1309));
   NAND2_X1 U791 (.A1(REGISTERS[202]),
	.A2(n4022),
	.ZN(n285));
   OAI21_X1 U792 (.A(n286),
	.B1(FE_OFN85_n4022),
	.B2(n60),
	.ZN(n1310));
   NAND2_X1 U793 (.A1(REGISTERS[203]),
	.A2(FE_OFN85_n4022),
	.ZN(n286));
   OAI21_X1 U794 (.A(n287),
	.B1(n4022),
	.B2(n62),
	.ZN(n1311));
   NAND2_X1 U795 (.A1(REGISTERS[204]),
	.A2(n4022),
	.ZN(n287));
   OAI21_X1 U796 (.A(n289),
	.B1(FE_OFN85_n4022),
	.B2(n66),
	.ZN(n1313));
   NAND2_X1 U797 (.A1(REGISTERS[206]),
	.A2(FE_OFN85_n4022),
	.ZN(n289));
   OAI21_X1 U798 (.A(n290),
	.B1(n4022),
	.B2(n68),
	.ZN(n1314));
   NAND2_X1 U799 (.A1(REGISTERS[207]),
	.A2(n4022),
	.ZN(n290));
   OAI21_X1 U800 (.A(n316),
	.B1(FE_OFN72_n4021),
	.B2(n52),
	.ZN(n1338));
   NAND2_X1 U801 (.A1(REGISTERS[231]),
	.A2(FE_OFN72_n4021),
	.ZN(n316));
   OAI21_X1 U802 (.A(n317),
	.B1(n4021),
	.B2(n54),
	.ZN(n1339));
   NAND2_X1 U803 (.A1(REGISTERS[232]),
	.A2(n4021),
	.ZN(n317));
   OAI21_X1 U804 (.A(n318),
	.B1(FE_OFN72_n4021),
	.B2(n56),
	.ZN(n1340));
   NAND2_X1 U805 (.A1(REGISTERS[233]),
	.A2(FE_OFN72_n4021),
	.ZN(n318));
   OAI21_X1 U806 (.A(n319),
	.B1(n4021),
	.B2(n58),
	.ZN(n1341));
   NAND2_X1 U807 (.A1(REGISTERS[234]),
	.A2(n4021),
	.ZN(n319));
   OAI21_X1 U808 (.A(n320),
	.B1(FE_OFN72_n4021),
	.B2(n60),
	.ZN(n1342));
   NAND2_X1 U809 (.A1(REGISTERS[235]),
	.A2(FE_OFN72_n4021),
	.ZN(n320));
   OAI21_X1 U810 (.A(n321),
	.B1(n4021),
	.B2(n62),
	.ZN(n1343));
   NAND2_X1 U811 (.A1(REGISTERS[236]),
	.A2(n4021),
	.ZN(n321));
   OAI21_X1 U812 (.A(n323),
	.B1(FE_OFN72_n4021),
	.B2(n66),
	.ZN(n1345));
   NAND2_X1 U813 (.A1(REGISTERS[238]),
	.A2(FE_OFN72_n4021),
	.ZN(n323));
   OAI21_X1 U814 (.A(n324),
	.B1(n4021),
	.B2(n68),
	.ZN(n1346));
   NAND2_X1 U815 (.A1(REGISTERS[239]),
	.A2(n4021),
	.ZN(n324));
   OAI21_X1 U816 (.A(n343),
	.B1(FE_OFN60_n4036),
	.B2(n38),
	.ZN(n1363));
   NAND2_X1 U817 (.A1(REGISTERS[256]),
	.A2(FE_OFN60_n4036),
	.ZN(n343));
   OAI21_X1 U818 (.A(n345),
	.B1(FE_OFN60_n4036),
	.B2(n42),
	.ZN(n1365));
   NAND2_X1 U819 (.A1(REGISTERS[258]),
	.A2(FE_OFN60_n4036),
	.ZN(n345));
   OAI21_X1 U820 (.A(n348),
	.B1(FE_OFN60_n4036),
	.B2(n48),
	.ZN(n1368));
   NAND2_X1 U821 (.A1(REGISTERS[261]),
	.A2(FE_OFN60_n4036),
	.ZN(n348));
   OAI21_X1 U822 (.A(n349),
	.B1(n4036),
	.B2(n50),
	.ZN(n1369));
   NAND2_X1 U823 (.A1(REGISTERS[262]),
	.A2(n4036),
	.ZN(n349));
   OAI21_X1 U824 (.A(n356),
	.B1(n4036),
	.B2(n64),
	.ZN(n1376));
   NAND2_X1 U825 (.A1(REGISTERS[269]),
	.A2(n4036),
	.ZN(n356));
   OAI21_X1 U826 (.A(n359),
	.B1(n4036),
	.B2(n70),
	.ZN(n1379));
   NAND2_X1 U827 (.A1(REGISTERS[272]),
	.A2(n4036),
	.ZN(n359));
   OAI21_X1 U828 (.A(n360),
	.B1(FE_OFN60_n4036),
	.B2(n72),
	.ZN(n1380));
   NAND2_X1 U829 (.A1(REGISTERS[273]),
	.A2(FE_OFN60_n4036),
	.ZN(n360));
   OAI21_X1 U830 (.A(n361),
	.B1(n4036),
	.B2(n74),
	.ZN(n1381));
   NAND2_X1 U831 (.A1(REGISTERS[274]),
	.A2(n4036),
	.ZN(n361));
   OAI21_X1 U832 (.A(n362),
	.B1(FE_OFN60_n4036),
	.B2(n76),
	.ZN(n1382));
   NAND2_X1 U833 (.A1(REGISTERS[275]),
	.A2(FE_OFN60_n4036),
	.ZN(n362));
   OAI21_X1 U834 (.A(n363),
	.B1(n4036),
	.B2(n78),
	.ZN(n1383));
   NAND2_X1 U835 (.A1(REGISTERS[276]),
	.A2(n4036),
	.ZN(n363));
   OAI21_X1 U836 (.A(n364),
	.B1(FE_OFN60_n4036),
	.B2(n80),
	.ZN(n1384));
   NAND2_X1 U837 (.A1(REGISTERS[277]),
	.A2(FE_OFN60_n4036),
	.ZN(n364));
   OAI21_X1 U838 (.A(n365),
	.B1(FE_OFN60_n4036),
	.B2(n82),
	.ZN(n1385));
   NAND2_X1 U839 (.A1(REGISTERS[278]),
	.A2(FE_OFN60_n4036),
	.ZN(n365));
   OAI21_X1 U840 (.A(n366),
	.B1(FE_OFN60_n4036),
	.B2(n84),
	.ZN(n1386));
   NAND2_X1 U841 (.A1(REGISTERS[279]),
	.A2(FE_OFN60_n4036),
	.ZN(n366));
   OAI21_X1 U842 (.A(n367),
	.B1(n4036),
	.B2(n86),
	.ZN(n1387));
   NAND2_X1 U843 (.A1(REGISTERS[280]),
	.A2(n4036),
	.ZN(n367));
   OAI21_X1 U844 (.A(n368),
	.B1(FE_OFN60_n4036),
	.B2(n88),
	.ZN(n1388));
   NAND2_X1 U845 (.A1(REGISTERS[281]),
	.A2(FE_OFN60_n4036),
	.ZN(n368));
   OAI21_X1 U846 (.A(n369),
	.B1(n4036),
	.B2(n90),
	.ZN(n1389));
   NAND2_X1 U847 (.A1(REGISTERS[282]),
	.A2(n4036),
	.ZN(n369));
   OAI21_X1 U848 (.A(n370),
	.B1(FE_OFN60_n4036),
	.B2(n92),
	.ZN(n1390));
   NAND2_X1 U849 (.A1(REGISTERS[283]),
	.A2(FE_OFN60_n4036),
	.ZN(n370));
   OAI21_X1 U850 (.A(n371),
	.B1(FE_OFN60_n4036),
	.B2(n94),
	.ZN(n1391));
   NAND2_X1 U851 (.A1(REGISTERS[284]),
	.A2(FE_OFN60_n4036),
	.ZN(n371));
   OAI21_X1 U852 (.A(n377),
	.B1(FE_OFN80_n4035),
	.B2(n38),
	.ZN(n1395));
   NAND2_X1 U853 (.A1(REGISTERS[288]),
	.A2(FE_OFN80_n4035),
	.ZN(n377));
   OAI21_X1 U854 (.A(n379),
	.B1(FE_OFN80_n4035),
	.B2(n42),
	.ZN(n1397));
   NAND2_X1 U855 (.A1(REGISTERS[290]),
	.A2(FE_OFN80_n4035),
	.ZN(n379));
   OAI21_X1 U856 (.A(n382),
	.B1(FE_OFN80_n4035),
	.B2(n48),
	.ZN(n1400));
   NAND2_X1 U857 (.A1(REGISTERS[293]),
	.A2(FE_OFN80_n4035),
	.ZN(n382));
   OAI21_X1 U858 (.A(n383),
	.B1(n4035),
	.B2(n50),
	.ZN(n1401));
   NAND2_X1 U859 (.A1(REGISTERS[294]),
	.A2(n4035),
	.ZN(n383));
   OAI21_X1 U860 (.A(n390),
	.B1(n4035),
	.B2(n64),
	.ZN(n1408));
   NAND2_X1 U861 (.A1(REGISTERS[301]),
	.A2(n4035),
	.ZN(n390));
   OAI21_X1 U862 (.A(n393),
	.B1(FE_OFN80_n4035),
	.B2(n70),
	.ZN(n1411));
   NAND2_X1 U863 (.A1(REGISTERS[304]),
	.A2(FE_OFN80_n4035),
	.ZN(n393));
   OAI21_X1 U864 (.A(n394),
	.B1(FE_OFN80_n4035),
	.B2(n72),
	.ZN(n1412));
   NAND2_X1 U865 (.A1(REGISTERS[305]),
	.A2(FE_OFN80_n4035),
	.ZN(n394));
   OAI21_X1 U866 (.A(n395),
	.B1(n4035),
	.B2(n74),
	.ZN(n1413));
   NAND2_X1 U867 (.A1(REGISTERS[306]),
	.A2(n4035),
	.ZN(n395));
   OAI21_X1 U868 (.A(n396),
	.B1(FE_OFN80_n4035),
	.B2(n76),
	.ZN(n1414));
   NAND2_X1 U869 (.A1(REGISTERS[307]),
	.A2(FE_OFN80_n4035),
	.ZN(n396));
   OAI21_X1 U870 (.A(n397),
	.B1(n4035),
	.B2(n78),
	.ZN(n1415));
   NAND2_X1 U871 (.A1(REGISTERS[308]),
	.A2(n4035),
	.ZN(n397));
   OAI21_X1 U872 (.A(n398),
	.B1(FE_OFN80_n4035),
	.B2(n80),
	.ZN(n1416));
   NAND2_X1 U873 (.A1(REGISTERS[309]),
	.A2(FE_OFN80_n4035),
	.ZN(n398));
   OAI21_X1 U874 (.A(n399),
	.B1(FE_OFN80_n4035),
	.B2(n82),
	.ZN(n1417));
   NAND2_X1 U875 (.A1(REGISTERS[310]),
	.A2(FE_OFN80_n4035),
	.ZN(n399));
   OAI21_X1 U876 (.A(n400),
	.B1(FE_OFN80_n4035),
	.B2(n84),
	.ZN(n1418));
   NAND2_X1 U877 (.A1(REGISTERS[311]),
	.A2(FE_OFN80_n4035),
	.ZN(n400));
   OAI21_X1 U878 (.A(n401),
	.B1(n4035),
	.B2(n86),
	.ZN(n1419));
   NAND2_X1 U879 (.A1(REGISTERS[312]),
	.A2(n4035),
	.ZN(n401));
   OAI21_X1 U880 (.A(n402),
	.B1(FE_OFN80_n4035),
	.B2(n88),
	.ZN(n1420));
   NAND2_X1 U881 (.A1(REGISTERS[313]),
	.A2(FE_OFN80_n4035),
	.ZN(n402));
   OAI21_X1 U882 (.A(n403),
	.B1(n4035),
	.B2(n90),
	.ZN(n1421));
   NAND2_X1 U883 (.A1(REGISTERS[314]),
	.A2(n4035),
	.ZN(n403));
   OAI21_X1 U884 (.A(n404),
	.B1(FE_OFN80_n4035),
	.B2(n92),
	.ZN(n1422));
   NAND2_X1 U885 (.A1(REGISTERS[315]),
	.A2(FE_OFN80_n4035),
	.ZN(n404));
   OAI21_X1 U886 (.A(n405),
	.B1(FE_OFN80_n4035),
	.B2(n94),
	.ZN(n1423));
   NAND2_X1 U887 (.A1(REGISTERS[316]),
	.A2(FE_OFN80_n4035),
	.ZN(n405));
   OAI21_X1 U888 (.A(n410),
	.B1(FE_OFN59_n4034),
	.B2(n38),
	.ZN(n1427));
   NAND2_X1 U889 (.A1(REGISTERS[320]),
	.A2(FE_OFN59_n4034),
	.ZN(n410));
   OAI21_X1 U890 (.A(n412),
	.B1(FE_OFN59_n4034),
	.B2(n42),
	.ZN(n1429));
   NAND2_X1 U891 (.A1(REGISTERS[322]),
	.A2(FE_OFN59_n4034),
	.ZN(n412));
   OAI21_X1 U892 (.A(n415),
	.B1(FE_OFN59_n4034),
	.B2(n48),
	.ZN(n1432));
   NAND2_X1 U893 (.A1(REGISTERS[325]),
	.A2(FE_OFN59_n4034),
	.ZN(n415));
   OAI21_X1 U894 (.A(n416),
	.B1(FE_OFN59_n4034),
	.B2(n50),
	.ZN(n1433));
   NAND2_X1 U895 (.A1(REGISTERS[326]),
	.A2(FE_OFN59_n4034),
	.ZN(n416));
   OAI21_X1 U896 (.A(n423),
	.B1(FE_OFN59_n4034),
	.B2(n64),
	.ZN(n1440));
   NAND2_X1 U897 (.A1(REGISTERS[333]),
	.A2(FE_OFN59_n4034),
	.ZN(n423));
   OAI21_X1 U898 (.A(n426),
	.B1(n4034),
	.B2(n70),
	.ZN(n1443));
   NAND2_X1 U899 (.A1(REGISTERS[336]),
	.A2(n4034),
	.ZN(n426));
   OAI21_X1 U900 (.A(n427),
	.B1(FE_OFN59_n4034),
	.B2(n72),
	.ZN(n1444));
   NAND2_X1 U901 (.A1(REGISTERS[337]),
	.A2(FE_OFN59_n4034),
	.ZN(n427));
   OAI21_X1 U902 (.A(n428),
	.B1(FE_OFN59_n4034),
	.B2(n74),
	.ZN(n1445));
   NAND2_X1 U903 (.A1(REGISTERS[338]),
	.A2(FE_OFN59_n4034),
	.ZN(n428));
   OAI21_X1 U904 (.A(n429),
	.B1(FE_OFN59_n4034),
	.B2(n76),
	.ZN(n1446));
   NAND2_X1 U905 (.A1(REGISTERS[339]),
	.A2(FE_OFN59_n4034),
	.ZN(n429));
   OAI21_X1 U906 (.A(n430),
	.B1(FE_OFN59_n4034),
	.B2(n78),
	.ZN(n1447));
   NAND2_X1 U907 (.A1(REGISTERS[340]),
	.A2(FE_OFN59_n4034),
	.ZN(n430));
   OAI21_X1 U908 (.A(n431),
	.B1(FE_OFN59_n4034),
	.B2(n80),
	.ZN(n1448));
   NAND2_X1 U909 (.A1(REGISTERS[341]),
	.A2(FE_OFN59_n4034),
	.ZN(n431));
   OAI21_X1 U910 (.A(n432),
	.B1(FE_OFN59_n4034),
	.B2(n82),
	.ZN(n1449));
   NAND2_X1 U911 (.A1(REGISTERS[342]),
	.A2(FE_OFN59_n4034),
	.ZN(n432));
   OAI21_X1 U912 (.A(n433),
	.B1(FE_OFN59_n4034),
	.B2(n84),
	.ZN(n1450));
   NAND2_X1 U913 (.A1(REGISTERS[343]),
	.A2(FE_OFN59_n4034),
	.ZN(n433));
   OAI21_X1 U914 (.A(n434),
	.B1(FE_OFN59_n4034),
	.B2(n86),
	.ZN(n1451));
   NAND2_X1 U915 (.A1(REGISTERS[344]),
	.A2(FE_OFN59_n4034),
	.ZN(n434));
   OAI21_X1 U916 (.A(n435),
	.B1(FE_OFN59_n4034),
	.B2(n88),
	.ZN(n1452));
   NAND2_X1 U917 (.A1(REGISTERS[345]),
	.A2(FE_OFN59_n4034),
	.ZN(n435));
   OAI21_X1 U918 (.A(n436),
	.B1(FE_OFN59_n4034),
	.B2(n90),
	.ZN(n1453));
   NAND2_X1 U919 (.A1(REGISTERS[346]),
	.A2(FE_OFN59_n4034),
	.ZN(n436));
   OAI21_X1 U920 (.A(n437),
	.B1(FE_OFN59_n4034),
	.B2(n92),
	.ZN(n1454));
   NAND2_X1 U921 (.A1(REGISTERS[347]),
	.A2(FE_OFN59_n4034),
	.ZN(n437));
   OAI21_X1 U922 (.A(n438),
	.B1(FE_OFN59_n4034),
	.B2(n94),
	.ZN(n1455));
   NAND2_X1 U923 (.A1(REGISTERS[348]),
	.A2(FE_OFN59_n4034),
	.ZN(n438));
   OAI21_X1 U924 (.A(n443),
	.B1(FE_OFN70_n4033),
	.B2(n38),
	.ZN(n1459));
   NAND2_X1 U925 (.A1(REGISTERS[352]),
	.A2(FE_OFN70_n4033),
	.ZN(n443));
   OAI21_X1 U926 (.A(n445),
	.B1(FE_OFN70_n4033),
	.B2(n42),
	.ZN(n1461));
   NAND2_X1 U927 (.A1(REGISTERS[354]),
	.A2(FE_OFN70_n4033),
	.ZN(n445));
   OAI21_X1 U928 (.A(n448),
	.B1(FE_OFN70_n4033),
	.B2(n48),
	.ZN(n1464));
   NAND2_X1 U929 (.A1(REGISTERS[357]),
	.A2(FE_OFN70_n4033),
	.ZN(n448));
   OAI21_X1 U930 (.A(n449),
	.B1(FE_OFN70_n4033),
	.B2(n50),
	.ZN(n1465));
   NAND2_X1 U931 (.A1(REGISTERS[358]),
	.A2(FE_OFN70_n4033),
	.ZN(n449));
   OAI21_X1 U932 (.A(n456),
	.B1(FE_OFN70_n4033),
	.B2(n64),
	.ZN(n1472));
   NAND2_X1 U933 (.A1(REGISTERS[365]),
	.A2(FE_OFN70_n4033),
	.ZN(n456));
   OAI21_X1 U934 (.A(n459),
	.B1(FE_OFN70_n4033),
	.B2(n70),
	.ZN(n1475));
   NAND2_X1 U935 (.A1(REGISTERS[368]),
	.A2(FE_OFN70_n4033),
	.ZN(n459));
   OAI21_X1 U936 (.A(n460),
	.B1(FE_OFN70_n4033),
	.B2(n72),
	.ZN(n1476));
   NAND2_X1 U937 (.A1(REGISTERS[369]),
	.A2(FE_OFN70_n4033),
	.ZN(n460));
   OAI21_X1 U938 (.A(n461),
	.B1(FE_OFN70_n4033),
	.B2(n74),
	.ZN(n1477));
   NAND2_X1 U939 (.A1(REGISTERS[370]),
	.A2(FE_OFN70_n4033),
	.ZN(n461));
   OAI21_X1 U940 (.A(n462),
	.B1(FE_OFN70_n4033),
	.B2(n76),
	.ZN(n1478));
   NAND2_X1 U941 (.A1(REGISTERS[371]),
	.A2(FE_OFN70_n4033),
	.ZN(n462));
   OAI21_X1 U942 (.A(n463),
	.B1(FE_OFN70_n4033),
	.B2(n78),
	.ZN(n1479));
   NAND2_X1 U943 (.A1(REGISTERS[372]),
	.A2(FE_OFN70_n4033),
	.ZN(n463));
   OAI21_X1 U944 (.A(n464),
	.B1(FE_OFN70_n4033),
	.B2(n80),
	.ZN(n1480));
   NAND2_X1 U945 (.A1(REGISTERS[373]),
	.A2(FE_OFN70_n4033),
	.ZN(n464));
   OAI21_X1 U946 (.A(n465),
	.B1(FE_OFN70_n4033),
	.B2(n82),
	.ZN(n1481));
   NAND2_X1 U947 (.A1(REGISTERS[374]),
	.A2(FE_OFN70_n4033),
	.ZN(n465));
   OAI21_X1 U948 (.A(n466),
	.B1(FE_OFN70_n4033),
	.B2(n84),
	.ZN(n1482));
   NAND2_X1 U949 (.A1(REGISTERS[375]),
	.A2(FE_OFN70_n4033),
	.ZN(n466));
   OAI21_X1 U950 (.A(n467),
	.B1(FE_OFN70_n4033),
	.B2(n86),
	.ZN(n1483));
   NAND2_X1 U951 (.A1(REGISTERS[376]),
	.A2(FE_OFN70_n4033),
	.ZN(n467));
   OAI21_X1 U952 (.A(n468),
	.B1(FE_OFN70_n4033),
	.B2(n88),
	.ZN(n1484));
   NAND2_X1 U953 (.A1(REGISTERS[377]),
	.A2(FE_OFN70_n4033),
	.ZN(n468));
   OAI21_X1 U954 (.A(n469),
	.B1(FE_OFN70_n4033),
	.B2(n90),
	.ZN(n1485));
   NAND2_X1 U955 (.A1(REGISTERS[378]),
	.A2(FE_OFN70_n4033),
	.ZN(n469));
   OAI21_X1 U956 (.A(n470),
	.B1(FE_OFN70_n4033),
	.B2(n92),
	.ZN(n1486));
   NAND2_X1 U957 (.A1(REGISTERS[379]),
	.A2(FE_OFN70_n4033),
	.ZN(n470));
   OAI21_X1 U958 (.A(n471),
	.B1(FE_OFN70_n4033),
	.B2(n94),
	.ZN(n1487));
   NAND2_X1 U959 (.A1(REGISTERS[380]),
	.A2(FE_OFN70_n4033),
	.ZN(n471));
   OAI21_X1 U960 (.A(n476),
	.B1(FE_OFN87_n4032),
	.B2(n38),
	.ZN(n1491));
   NAND2_X1 U961 (.A1(REGISTERS[384]),
	.A2(FE_OFN87_n4032),
	.ZN(n476));
   OAI21_X1 U962 (.A(n478),
	.B1(FE_OFN87_n4032),
	.B2(n42),
	.ZN(n1493));
   NAND2_X1 U963 (.A1(REGISTERS[386]),
	.A2(FE_OFN87_n4032),
	.ZN(n478));
   OAI21_X1 U964 (.A(n481),
	.B1(FE_OFN87_n4032),
	.B2(n48),
	.ZN(n1496));
   NAND2_X1 U965 (.A1(REGISTERS[389]),
	.A2(FE_OFN87_n4032),
	.ZN(n481));
   OAI21_X1 U966 (.A(n482),
	.B1(n4032),
	.B2(n50),
	.ZN(n1497));
   NAND2_X1 U967 (.A1(REGISTERS[390]),
	.A2(n4032),
	.ZN(n482));
   OAI21_X1 U968 (.A(n489),
	.B1(n4032),
	.B2(n64),
	.ZN(n1504));
   NAND2_X1 U969 (.A1(REGISTERS[397]),
	.A2(n4032),
	.ZN(n489));
   OAI21_X1 U970 (.A(n492),
	.B1(FE_OFN87_n4032),
	.B2(n70),
	.ZN(n1507));
   NAND2_X1 U971 (.A1(REGISTERS[400]),
	.A2(FE_OFN87_n4032),
	.ZN(n492));
   OAI21_X1 U972 (.A(n493),
	.B1(FE_OFN87_n4032),
	.B2(n72),
	.ZN(n1508));
   NAND2_X1 U973 (.A1(REGISTERS[401]),
	.A2(FE_OFN87_n4032),
	.ZN(n493));
   OAI21_X1 U974 (.A(n494),
	.B1(n4032),
	.B2(n74),
	.ZN(n1509));
   NAND2_X1 U975 (.A1(REGISTERS[402]),
	.A2(n4032),
	.ZN(n494));
   OAI21_X1 U976 (.A(n495),
	.B1(FE_OFN87_n4032),
	.B2(n76),
	.ZN(n1510));
   NAND2_X1 U977 (.A1(REGISTERS[403]),
	.A2(FE_OFN87_n4032),
	.ZN(n495));
   OAI21_X1 U978 (.A(n496),
	.B1(n4032),
	.B2(n78),
	.ZN(n1511));
   NAND2_X1 U979 (.A1(REGISTERS[404]),
	.A2(n4032),
	.ZN(n496));
   OAI21_X1 U980 (.A(n497),
	.B1(FE_OFN87_n4032),
	.B2(n80),
	.ZN(n1512));
   NAND2_X1 U981 (.A1(REGISTERS[405]),
	.A2(FE_OFN87_n4032),
	.ZN(n497));
   OAI21_X1 U982 (.A(n498),
	.B1(FE_OFN87_n4032),
	.B2(n82),
	.ZN(n1513));
   NAND2_X1 U983 (.A1(REGISTERS[406]),
	.A2(FE_OFN87_n4032),
	.ZN(n498));
   OAI21_X1 U984 (.A(n499),
	.B1(FE_OFN87_n4032),
	.B2(n84),
	.ZN(n1514));
   NAND2_X1 U985 (.A1(REGISTERS[407]),
	.A2(FE_OFN87_n4032),
	.ZN(n499));
   OAI21_X1 U986 (.A(n500),
	.B1(n4032),
	.B2(n86),
	.ZN(n1515));
   NAND2_X1 U987 (.A1(REGISTERS[408]),
	.A2(n4032),
	.ZN(n500));
   OAI21_X1 U988 (.A(n501),
	.B1(FE_OFN87_n4032),
	.B2(n88),
	.ZN(n1516));
   NAND2_X1 U989 (.A1(REGISTERS[409]),
	.A2(FE_OFN87_n4032),
	.ZN(n501));
   OAI21_X1 U990 (.A(n502),
	.B1(n4032),
	.B2(n90),
	.ZN(n1517));
   NAND2_X1 U991 (.A1(REGISTERS[410]),
	.A2(n4032),
	.ZN(n502));
   OAI21_X1 U992 (.A(n503),
	.B1(FE_OFN87_n4032),
	.B2(n92),
	.ZN(n1518));
   NAND2_X1 U993 (.A1(REGISTERS[411]),
	.A2(FE_OFN87_n4032),
	.ZN(n503));
   OAI21_X1 U994 (.A(n504),
	.B1(FE_OFN87_n4032),
	.B2(n94),
	.ZN(n1519));
   NAND2_X1 U995 (.A1(REGISTERS[412]),
	.A2(FE_OFN87_n4032),
	.ZN(n504));
   OAI21_X1 U996 (.A(n509),
	.B1(FE_OFN63_n4031),
	.B2(n38),
	.ZN(n1523));
   NAND2_X1 U997 (.A1(REGISTERS[416]),
	.A2(FE_OFN63_n4031),
	.ZN(n509));
   OAI21_X1 U998 (.A(n511),
	.B1(FE_OFN63_n4031),
	.B2(n42),
	.ZN(n1525));
   NAND2_X1 U999 (.A1(REGISTERS[418]),
	.A2(FE_OFN63_n4031),
	.ZN(n511));
   OAI21_X1 U1000 (.A(n514),
	.B1(FE_OFN63_n4031),
	.B2(n48),
	.ZN(n1528));
   NAND2_X1 U1001 (.A1(REGISTERS[421]),
	.A2(FE_OFN63_n4031),
	.ZN(n514));
   OAI21_X1 U1002 (.A(n515),
	.B1(FE_OFN63_n4031),
	.B2(n50),
	.ZN(n1529));
   NAND2_X1 U1003 (.A1(REGISTERS[422]),
	.A2(FE_OFN63_n4031),
	.ZN(n515));
   OAI21_X1 U1004 (.A(n522),
	.B1(FE_OFN63_n4031),
	.B2(n64),
	.ZN(n1536));
   NAND2_X1 U1005 (.A1(REGISTERS[429]),
	.A2(FE_OFN63_n4031),
	.ZN(n522));
   OAI21_X1 U1006 (.A(n525),
	.B1(n4031),
	.B2(n70),
	.ZN(n1539));
   NAND2_X1 U1007 (.A1(REGISTERS[432]),
	.A2(n4031),
	.ZN(n525));
   OAI21_X1 U1008 (.A(n526),
	.B1(FE_OFN63_n4031),
	.B2(n72),
	.ZN(n1540));
   NAND2_X1 U1009 (.A1(REGISTERS[433]),
	.A2(FE_OFN63_n4031),
	.ZN(n526));
   OAI21_X1 U1010 (.A(n527),
	.B1(FE_OFN63_n4031),
	.B2(n74),
	.ZN(n1541));
   NAND2_X1 U1011 (.A1(REGISTERS[434]),
	.A2(FE_OFN63_n4031),
	.ZN(n527));
   OAI21_X1 U1012 (.A(n528),
	.B1(FE_OFN63_n4031),
	.B2(n76),
	.ZN(n1542));
   NAND2_X1 U1013 (.A1(REGISTERS[435]),
	.A2(FE_OFN63_n4031),
	.ZN(n528));
   OAI21_X1 U1014 (.A(n529),
	.B1(FE_OFN63_n4031),
	.B2(n78),
	.ZN(n1543));
   NAND2_X1 U1015 (.A1(REGISTERS[436]),
	.A2(FE_OFN63_n4031),
	.ZN(n529));
   OAI21_X1 U1016 (.A(n530),
	.B1(FE_OFN63_n4031),
	.B2(n80),
	.ZN(n1544));
   NAND2_X1 U1017 (.A1(REGISTERS[437]),
	.A2(FE_OFN63_n4031),
	.ZN(n530));
   OAI21_X1 U1018 (.A(n531),
	.B1(FE_OFN63_n4031),
	.B2(n82),
	.ZN(n1545));
   NAND2_X1 U1019 (.A1(REGISTERS[438]),
	.A2(FE_OFN63_n4031),
	.ZN(n531));
   OAI21_X1 U1020 (.A(n532),
	.B1(FE_OFN63_n4031),
	.B2(n84),
	.ZN(n1546));
   NAND2_X1 U1021 (.A1(REGISTERS[439]),
	.A2(FE_OFN63_n4031),
	.ZN(n532));
   OAI21_X1 U1022 (.A(n533),
	.B1(FE_OFN63_n4031),
	.B2(n86),
	.ZN(n1547));
   NAND2_X1 U1023 (.A1(REGISTERS[440]),
	.A2(FE_OFN63_n4031),
	.ZN(n533));
   OAI21_X1 U1024 (.A(n534),
	.B1(FE_OFN63_n4031),
	.B2(n88),
	.ZN(n1548));
   NAND2_X1 U1025 (.A1(REGISTERS[441]),
	.A2(FE_OFN63_n4031),
	.ZN(n534));
   OAI21_X1 U1026 (.A(n535),
	.B1(FE_OFN63_n4031),
	.B2(n90),
	.ZN(n1549));
   NAND2_X1 U1027 (.A1(REGISTERS[442]),
	.A2(FE_OFN63_n4031),
	.ZN(n535));
   OAI21_X1 U1028 (.A(n536),
	.B1(FE_OFN63_n4031),
	.B2(n92),
	.ZN(n1550));
   NAND2_X1 U1029 (.A1(REGISTERS[443]),
	.A2(FE_OFN63_n4031),
	.ZN(n536));
   OAI21_X1 U1030 (.A(n537),
	.B1(FE_OFN63_n4031),
	.B2(n94),
	.ZN(n1551));
   NAND2_X1 U1031 (.A1(REGISTERS[444]),
	.A2(FE_OFN63_n4031),
	.ZN(n537));
   OAI21_X1 U1032 (.A(n542),
	.B1(FE_OFN81_n4030),
	.B2(n38),
	.ZN(n1555));
   NAND2_X1 U1033 (.A1(REGISTERS[448]),
	.A2(FE_OFN81_n4030),
	.ZN(n542));
   OAI21_X1 U1034 (.A(n544),
	.B1(FE_OFN81_n4030),
	.B2(n42),
	.ZN(n1557));
   NAND2_X1 U1035 (.A1(REGISTERS[450]),
	.A2(FE_OFN81_n4030),
	.ZN(n544));
   OAI21_X1 U1036 (.A(n547),
	.B1(FE_OFN81_n4030),
	.B2(n48),
	.ZN(n1560));
   NAND2_X1 U1037 (.A1(REGISTERS[453]),
	.A2(FE_OFN81_n4030),
	.ZN(n547));
   OAI21_X1 U1038 (.A(n548),
	.B1(n4030),
	.B2(n50),
	.ZN(n1561));
   NAND2_X1 U1039 (.A1(REGISTERS[454]),
	.A2(n4030),
	.ZN(n548));
   OAI21_X1 U1040 (.A(n555),
	.B1(n4030),
	.B2(n64),
	.ZN(n1568));
   NAND2_X1 U1041 (.A1(REGISTERS[461]),
	.A2(n4030),
	.ZN(n555));
   OAI21_X1 U1042 (.A(n558),
	.B1(FE_OFN81_n4030),
	.B2(n70),
	.ZN(n1571));
   NAND2_X1 U1043 (.A1(REGISTERS[464]),
	.A2(FE_OFN81_n4030),
	.ZN(n558));
   OAI21_X1 U1044 (.A(n559),
	.B1(FE_OFN81_n4030),
	.B2(n72),
	.ZN(n1572));
   NAND2_X1 U1045 (.A1(REGISTERS[465]),
	.A2(FE_OFN81_n4030),
	.ZN(n559));
   OAI21_X1 U1046 (.A(n560),
	.B1(n4030),
	.B2(n74),
	.ZN(n1573));
   NAND2_X1 U1047 (.A1(REGISTERS[466]),
	.A2(n4030),
	.ZN(n560));
   OAI21_X1 U1048 (.A(n561),
	.B1(FE_OFN81_n4030),
	.B2(n76),
	.ZN(n1574));
   NAND2_X1 U1049 (.A1(REGISTERS[467]),
	.A2(FE_OFN81_n4030),
	.ZN(n561));
   OAI21_X1 U1050 (.A(n562),
	.B1(n4030),
	.B2(n78),
	.ZN(n1575));
   NAND2_X1 U1051 (.A1(REGISTERS[468]),
	.A2(n4030),
	.ZN(n562));
   OAI21_X1 U1052 (.A(n563),
	.B1(FE_OFN81_n4030),
	.B2(n80),
	.ZN(n1576));
   NAND2_X1 U1053 (.A1(REGISTERS[469]),
	.A2(FE_OFN81_n4030),
	.ZN(n563));
   OAI21_X1 U1054 (.A(n564),
	.B1(FE_OFN81_n4030),
	.B2(n82),
	.ZN(n1577));
   NAND2_X1 U1055 (.A1(REGISTERS[470]),
	.A2(FE_OFN81_n4030),
	.ZN(n564));
   OAI21_X1 U1056 (.A(n565),
	.B1(FE_OFN81_n4030),
	.B2(n84),
	.ZN(n1578));
   NAND2_X1 U1057 (.A1(REGISTERS[471]),
	.A2(FE_OFN81_n4030),
	.ZN(n565));
   OAI21_X1 U1058 (.A(n566),
	.B1(n4030),
	.B2(n86),
	.ZN(n1579));
   NAND2_X1 U1059 (.A1(REGISTERS[472]),
	.A2(n4030),
	.ZN(n566));
   OAI21_X1 U1060 (.A(n567),
	.B1(FE_OFN81_n4030),
	.B2(n88),
	.ZN(n1580));
   NAND2_X1 U1061 (.A1(REGISTERS[473]),
	.A2(FE_OFN81_n4030),
	.ZN(n567));
   OAI21_X1 U1062 (.A(n568),
	.B1(n4030),
	.B2(n90),
	.ZN(n1581));
   NAND2_X1 U1063 (.A1(REGISTERS[474]),
	.A2(n4030),
	.ZN(n568));
   OAI21_X1 U1064 (.A(n569),
	.B1(FE_OFN81_n4030),
	.B2(n92),
	.ZN(n1582));
   NAND2_X1 U1065 (.A1(REGISTERS[475]),
	.A2(FE_OFN81_n4030),
	.ZN(n569));
   OAI21_X1 U1066 (.A(n570),
	.B1(FE_OFN81_n4030),
	.B2(n94),
	.ZN(n1583));
   NAND2_X1 U1067 (.A1(REGISTERS[476]),
	.A2(FE_OFN81_n4030),
	.ZN(n570));
   OAI21_X1 U1068 (.A(n575),
	.B1(n4029),
	.B2(n38),
	.ZN(n1587));
   NAND2_X1 U1069 (.A1(REGISTERS[480]),
	.A2(n4029),
	.ZN(n575));
   OAI21_X1 U1070 (.A(n577),
	.B1(FE_OFN67_n4029),
	.B2(n42),
	.ZN(n1589));
   NAND2_X1 U1071 (.A1(REGISTERS[482]),
	.A2(FE_OFN67_n4029),
	.ZN(n577));
   OAI21_X1 U1072 (.A(n580),
	.B1(FE_OFN67_n4029),
	.B2(n48),
	.ZN(n1592));
   NAND2_X1 U1073 (.A1(REGISTERS[485]),
	.A2(FE_OFN67_n4029),
	.ZN(n580));
   OAI21_X1 U1074 (.A(n581),
	.B1(n4029),
	.B2(n50),
	.ZN(n1593));
   NAND2_X1 U1075 (.A1(REGISTERS[486]),
	.A2(n4029),
	.ZN(n581));
   OAI21_X1 U1076 (.A(n588),
	.B1(n4029),
	.B2(n64),
	.ZN(n1600));
   NAND2_X1 U1077 (.A1(REGISTERS[493]),
	.A2(n4029),
	.ZN(n588));
   OAI21_X1 U1078 (.A(n591),
	.B1(FE_OFN67_n4029),
	.B2(n70),
	.ZN(n1603));
   NAND2_X1 U1079 (.A1(REGISTERS[496]),
	.A2(FE_OFN67_n4029),
	.ZN(n591));
   OAI21_X1 U1080 (.A(n592),
	.B1(FE_OFN67_n4029),
	.B2(n72),
	.ZN(n1604));
   NAND2_X1 U1081 (.A1(REGISTERS[497]),
	.A2(FE_OFN67_n4029),
	.ZN(n592));
   OAI21_X1 U1082 (.A(n593),
	.B1(n4029),
	.B2(n74),
	.ZN(n1605));
   NAND2_X1 U1083 (.A1(REGISTERS[498]),
	.A2(n4029),
	.ZN(n593));
   OAI21_X1 U1084 (.A(n594),
	.B1(FE_OFN67_n4029),
	.B2(n76),
	.ZN(n1606));
   NAND2_X1 U1085 (.A1(REGISTERS[499]),
	.A2(FE_OFN67_n4029),
	.ZN(n594));
   OAI21_X1 U1086 (.A(n595),
	.B1(n4029),
	.B2(n78),
	.ZN(n1607));
   NAND2_X1 U1087 (.A1(REGISTERS[500]),
	.A2(n4029),
	.ZN(n595));
   OAI21_X1 U1088 (.A(n596),
	.B1(FE_OFN67_n4029),
	.B2(n80),
	.ZN(n1608));
   NAND2_X1 U1089 (.A1(REGISTERS[501]),
	.A2(FE_OFN67_n4029),
	.ZN(n596));
   OAI21_X1 U1090 (.A(n597),
	.B1(FE_OFN67_n4029),
	.B2(n82),
	.ZN(n1609));
   NAND2_X1 U1091 (.A1(REGISTERS[502]),
	.A2(FE_OFN67_n4029),
	.ZN(n597));
   OAI21_X1 U1092 (.A(n598),
	.B1(FE_OFN67_n4029),
	.B2(n84),
	.ZN(n1610));
   NAND2_X1 U1093 (.A1(REGISTERS[503]),
	.A2(FE_OFN67_n4029),
	.ZN(n598));
   OAI21_X1 U1094 (.A(n599),
	.B1(n4029),
	.B2(n86),
	.ZN(n1611));
   NAND2_X1 U1095 (.A1(REGISTERS[504]),
	.A2(n4029),
	.ZN(n599));
   OAI21_X1 U1096 (.A(n600),
	.B1(FE_OFN67_n4029),
	.B2(n88),
	.ZN(n1612));
   NAND2_X1 U1097 (.A1(REGISTERS[505]),
	.A2(FE_OFN67_n4029),
	.ZN(n600));
   OAI21_X1 U1098 (.A(n601),
	.B1(n4029),
	.B2(n90),
	.ZN(n1613));
   NAND2_X1 U1099 (.A1(REGISTERS[506]),
	.A2(n4029),
	.ZN(n601));
   OAI21_X1 U1100 (.A(n602),
	.B1(FE_OFN67_n4029),
	.B2(n92),
	.ZN(n1614));
   NAND2_X1 U1101 (.A1(REGISTERS[507]),
	.A2(FE_OFN67_n4029),
	.ZN(n602));
   OAI21_X1 U1102 (.A(n603),
	.B1(FE_OFN67_n4029),
	.B2(n94),
	.ZN(n1615));
   NAND2_X1 U1103 (.A1(REGISTERS[508]),
	.A2(FE_OFN67_n4029),
	.ZN(n603));
   OAI21_X1 U1104 (.A(n608),
	.B1(n4019),
	.B2(n38),
	.ZN(n1619));
   NAND2_X1 U1105 (.A1(REGISTERS[512]),
	.A2(n4019),
	.ZN(n608));
   OAI21_X1 U1106 (.A(n610),
	.B1(FE_OFN61_n4019),
	.B2(n42),
	.ZN(n1621));
   NAND2_X1 U1107 (.A1(REGISTERS[514]),
	.A2(FE_OFN61_n4019),
	.ZN(n610));
   OAI21_X1 U1108 (.A(n613),
	.B1(FE_OFN61_n4019),
	.B2(n48),
	.ZN(n1624));
   NAND2_X1 U1109 (.A1(REGISTERS[517]),
	.A2(FE_OFN61_n4019),
	.ZN(n613));
   OAI21_X1 U1110 (.A(n614),
	.B1(n4019),
	.B2(n50),
	.ZN(n1625));
   NAND2_X1 U1111 (.A1(REGISTERS[518]),
	.A2(n4019),
	.ZN(n614));
   OAI21_X1 U1112 (.A(n621),
	.B1(n4019),
	.B2(n64),
	.ZN(n1632));
   NAND2_X1 U1113 (.A1(REGISTERS[525]),
	.A2(n4019),
	.ZN(n621));
   OAI21_X1 U1114 (.A(n624),
	.B1(n4019),
	.B2(n70),
	.ZN(n1635));
   NAND2_X1 U1115 (.A1(REGISTERS[528]),
	.A2(FE_OFN61_n4019),
	.ZN(n624));
   OAI21_X1 U1116 (.A(n625),
	.B1(FE_OFN61_n4019),
	.B2(n72),
	.ZN(n1636));
   NAND2_X1 U1117 (.A1(REGISTERS[529]),
	.A2(FE_OFN61_n4019),
	.ZN(n625));
   OAI21_X1 U1118 (.A(n626),
	.B1(n4019),
	.B2(n74),
	.ZN(n1637));
   NAND2_X1 U1119 (.A1(REGISTERS[530]),
	.A2(n4019),
	.ZN(n626));
   OAI21_X1 U1120 (.A(n627),
	.B1(FE_OFN61_n4019),
	.B2(n76),
	.ZN(n1638));
   NAND2_X1 U1121 (.A1(REGISTERS[531]),
	.A2(FE_OFN61_n4019),
	.ZN(n627));
   OAI21_X1 U1122 (.A(n628),
	.B1(FE_OFN61_n4019),
	.B2(n78),
	.ZN(n1639));
   NAND2_X1 U1123 (.A1(REGISTERS[532]),
	.A2(FE_OFN61_n4019),
	.ZN(n628));
   OAI21_X1 U1124 (.A(n629),
	.B1(FE_OFN61_n4019),
	.B2(n80),
	.ZN(n1640));
   NAND2_X1 U1125 (.A1(REGISTERS[533]),
	.A2(FE_OFN61_n4019),
	.ZN(n629));
   OAI21_X1 U1126 (.A(n630),
	.B1(FE_OFN61_n4019),
	.B2(n82),
	.ZN(n1641));
   NAND2_X1 U1127 (.A1(REGISTERS[534]),
	.A2(FE_OFN61_n4019),
	.ZN(n630));
   OAI21_X1 U1128 (.A(n631),
	.B1(FE_OFN61_n4019),
	.B2(n84),
	.ZN(n1642));
   NAND2_X1 U1129 (.A1(REGISTERS[535]),
	.A2(FE_OFN61_n4019),
	.ZN(n631));
   OAI21_X1 U1130 (.A(n632),
	.B1(FE_OFN61_n4019),
	.B2(n86),
	.ZN(n1643));
   NAND2_X1 U1131 (.A1(REGISTERS[536]),
	.A2(FE_OFN61_n4019),
	.ZN(n632));
   OAI21_X1 U1132 (.A(n633),
	.B1(FE_OFN61_n4019),
	.B2(n88),
	.ZN(n1644));
   NAND2_X1 U1133 (.A1(REGISTERS[537]),
	.A2(FE_OFN61_n4019),
	.ZN(n633));
   OAI21_X1 U1134 (.A(n634),
	.B1(FE_OFN61_n4019),
	.B2(n90),
	.ZN(n1645));
   NAND2_X1 U1135 (.A1(REGISTERS[538]),
	.A2(FE_OFN61_n4019),
	.ZN(n634));
   OAI21_X1 U1136 (.A(n635),
	.B1(FE_OFN61_n4019),
	.B2(n92),
	.ZN(n1646));
   NAND2_X1 U1137 (.A1(REGISTERS[539]),
	.A2(FE_OFN61_n4019),
	.ZN(n635));
   OAI21_X1 U1138 (.A(n636),
	.B1(FE_OFN61_n4019),
	.B2(n94),
	.ZN(n1647));
   NAND2_X1 U1139 (.A1(REGISTERS[540]),
	.A2(FE_OFN61_n4019),
	.ZN(n636));
   OAI21_X1 U1140 (.A(n642),
	.B1(FE_OFN65_n4018),
	.B2(n38),
	.ZN(n1651));
   NAND2_X1 U1141 (.A1(REGISTERS[544]),
	.A2(FE_OFN65_n4018),
	.ZN(n642));
   OAI21_X1 U1142 (.A(n644),
	.B1(FE_OFN65_n4018),
	.B2(n42),
	.ZN(n1653));
   NAND2_X1 U1143 (.A1(REGISTERS[546]),
	.A2(FE_OFN65_n4018),
	.ZN(n644));
   OAI21_X1 U1144 (.A(n647),
	.B1(n4018),
	.B2(n48),
	.ZN(n1656));
   NAND2_X1 U1145 (.A1(REGISTERS[549]),
	.A2(n4018),
	.ZN(n647));
   OAI21_X1 U1146 (.A(n648),
	.B1(FE_OFN65_n4018),
	.B2(n50),
	.ZN(n1657));
   NAND2_X1 U1147 (.A1(REGISTERS[550]),
	.A2(FE_OFN65_n4018),
	.ZN(n648));
   OAI21_X1 U1148 (.A(n655),
	.B1(FE_OFN65_n4018),
	.B2(n64),
	.ZN(n1664));
   NAND2_X1 U1149 (.A1(REGISTERS[557]),
	.A2(FE_OFN65_n4018),
	.ZN(n655));
   OAI21_X1 U1150 (.A(n658),
	.B1(n4018),
	.B2(n70),
	.ZN(n1667));
   NAND2_X1 U1151 (.A1(REGISTERS[560]),
	.A2(n4018),
	.ZN(n658));
   OAI21_X1 U1152 (.A(n659),
	.B1(FE_OFN65_n4018),
	.B2(n72),
	.ZN(n1668));
   NAND2_X1 U1153 (.A1(REGISTERS[561]),
	.A2(FE_OFN65_n4018),
	.ZN(n659));
   OAI21_X1 U1154 (.A(n660),
	.B1(FE_OFN65_n4018),
	.B2(n74),
	.ZN(n1669));
   NAND2_X1 U1155 (.A1(REGISTERS[562]),
	.A2(FE_OFN65_n4018),
	.ZN(n660));
   OAI21_X1 U1156 (.A(n661),
	.B1(FE_OFN65_n4018),
	.B2(n76),
	.ZN(n1670));
   NAND2_X1 U1157 (.A1(REGISTERS[563]),
	.A2(FE_OFN65_n4018),
	.ZN(n661));
   OAI21_X1 U1158 (.A(n662),
	.B1(FE_OFN65_n4018),
	.B2(n78),
	.ZN(n1671));
   NAND2_X1 U1159 (.A1(REGISTERS[564]),
	.A2(FE_OFN65_n4018),
	.ZN(n662));
   OAI21_X1 U1160 (.A(n663),
	.B1(FE_OFN65_n4018),
	.B2(n80),
	.ZN(n1672));
   NAND2_X1 U1161 (.A1(REGISTERS[565]),
	.A2(FE_OFN65_n4018),
	.ZN(n663));
   OAI21_X1 U1162 (.A(n664),
	.B1(FE_OFN65_n4018),
	.B2(n82),
	.ZN(n1673));
   NAND2_X1 U1163 (.A1(REGISTERS[566]),
	.A2(FE_OFN65_n4018),
	.ZN(n664));
   OAI21_X1 U1164 (.A(n665),
	.B1(FE_OFN65_n4018),
	.B2(n84),
	.ZN(n1674));
   NAND2_X1 U1165 (.A1(REGISTERS[567]),
	.A2(FE_OFN65_n4018),
	.ZN(n665));
   OAI21_X1 U1166 (.A(n666),
	.B1(FE_OFN65_n4018),
	.B2(n86),
	.ZN(n1675));
   NAND2_X1 U1167 (.A1(REGISTERS[568]),
	.A2(FE_OFN65_n4018),
	.ZN(n666));
   OAI21_X1 U1168 (.A(n667),
	.B1(FE_OFN65_n4018),
	.B2(n88),
	.ZN(n1676));
   NAND2_X1 U1169 (.A1(REGISTERS[569]),
	.A2(FE_OFN65_n4018),
	.ZN(n667));
   OAI21_X1 U1170 (.A(n668),
	.B1(FE_OFN65_n4018),
	.B2(n90),
	.ZN(n1677));
   NAND2_X1 U1171 (.A1(REGISTERS[570]),
	.A2(FE_OFN65_n4018),
	.ZN(n668));
   OAI21_X1 U1172 (.A(n669),
	.B1(FE_OFN65_n4018),
	.B2(n92),
	.ZN(n1678));
   NAND2_X1 U1173 (.A1(REGISTERS[571]),
	.A2(FE_OFN65_n4018),
	.ZN(n669));
   OAI21_X1 U1174 (.A(n670),
	.B1(FE_OFN65_n4018),
	.B2(n94),
	.ZN(n1679));
   NAND2_X1 U1175 (.A1(REGISTERS[572]),
	.A2(FE_OFN65_n4018),
	.ZN(n670));
   OAI21_X1 U1176 (.A(n675),
	.B1(n4017),
	.B2(n38),
	.ZN(n1683));
   NAND2_X1 U1177 (.A1(REGISTERS[576]),
	.A2(n4017),
	.ZN(n675));
   OAI21_X1 U1178 (.A(n677),
	.B1(FE_OFN66_n4017),
	.B2(n42),
	.ZN(n1685));
   NAND2_X1 U1179 (.A1(REGISTERS[578]),
	.A2(FE_OFN66_n4017),
	.ZN(n677));
   OAI21_X1 U1180 (.A(n680),
	.B1(FE_OFN66_n4017),
	.B2(n48),
	.ZN(n1688));
   NAND2_X1 U1181 (.A1(REGISTERS[581]),
	.A2(FE_OFN66_n4017),
	.ZN(n680));
   OAI21_X1 U1182 (.A(n681),
	.B1(n4017),
	.B2(n50),
	.ZN(n1689));
   NAND2_X1 U1183 (.A1(REGISTERS[582]),
	.A2(n4017),
	.ZN(n681));
   OAI21_X1 U1184 (.A(n688),
	.B1(n4017),
	.B2(n64),
	.ZN(n1696));
   NAND2_X1 U1185 (.A1(REGISTERS[589]),
	.A2(n4017),
	.ZN(n688));
   OAI21_X1 U1186 (.A(n691),
	.B1(FE_OFN66_n4017),
	.B2(n70),
	.ZN(n1699));
   NAND2_X1 U1187 (.A1(REGISTERS[592]),
	.A2(FE_OFN66_n4017),
	.ZN(n691));
   OAI21_X1 U1188 (.A(n692),
	.B1(FE_OFN66_n4017),
	.B2(n72),
	.ZN(n1700));
   NAND2_X1 U1189 (.A1(REGISTERS[593]),
	.A2(FE_OFN66_n4017),
	.ZN(n692));
   OAI21_X1 U1190 (.A(n693),
	.B1(n4017),
	.B2(n74),
	.ZN(n1701));
   NAND2_X1 U1191 (.A1(REGISTERS[594]),
	.A2(n4017),
	.ZN(n693));
   OAI21_X1 U1192 (.A(n694),
	.B1(FE_OFN66_n4017),
	.B2(n76),
	.ZN(n1702));
   NAND2_X1 U1193 (.A1(REGISTERS[595]),
	.A2(FE_OFN66_n4017),
	.ZN(n694));
   OAI21_X1 U1194 (.A(n695),
	.B1(FE_OFN66_n4017),
	.B2(n78),
	.ZN(n1703));
   NAND2_X1 U1195 (.A1(REGISTERS[596]),
	.A2(FE_OFN66_n4017),
	.ZN(n695));
   OAI21_X1 U1196 (.A(n696),
	.B1(FE_OFN66_n4017),
	.B2(n80),
	.ZN(n1704));
   NAND2_X1 U1197 (.A1(REGISTERS[597]),
	.A2(FE_OFN66_n4017),
	.ZN(n696));
   OAI21_X1 U1198 (.A(n697),
	.B1(FE_OFN66_n4017),
	.B2(n82),
	.ZN(n1705));
   NAND2_X1 U1199 (.A1(REGISTERS[598]),
	.A2(FE_OFN66_n4017),
	.ZN(n697));
   OAI21_X1 U1200 (.A(n698),
	.B1(FE_OFN66_n4017),
	.B2(n84),
	.ZN(n1706));
   NAND2_X1 U1201 (.A1(REGISTERS[599]),
	.A2(FE_OFN66_n4017),
	.ZN(n698));
   OAI21_X1 U1202 (.A(n699),
	.B1(FE_OFN66_n4017),
	.B2(n86),
	.ZN(n1707));
   NAND2_X1 U1203 (.A1(REGISTERS[600]),
	.A2(FE_OFN66_n4017),
	.ZN(n699));
   OAI21_X1 U1204 (.A(n700),
	.B1(FE_OFN66_n4017),
	.B2(n88),
	.ZN(n1708));
   NAND2_X1 U1205 (.A1(REGISTERS[601]),
	.A2(FE_OFN66_n4017),
	.ZN(n700));
   OAI21_X1 U1206 (.A(n701),
	.B1(FE_OFN66_n4017),
	.B2(n90),
	.ZN(n1709));
   NAND2_X1 U1207 (.A1(REGISTERS[602]),
	.A2(FE_OFN66_n4017),
	.ZN(n701));
   OAI21_X1 U1208 (.A(n702),
	.B1(FE_OFN66_n4017),
	.B2(n92),
	.ZN(n1710));
   NAND2_X1 U1209 (.A1(REGISTERS[603]),
	.A2(FE_OFN66_n4017),
	.ZN(n702));
   OAI21_X1 U1210 (.A(n703),
	.B1(FE_OFN66_n4017),
	.B2(n94),
	.ZN(n1711));
   NAND2_X1 U1211 (.A1(REGISTERS[604]),
	.A2(FE_OFN66_n4017),
	.ZN(n703));
   OAI21_X1 U1212 (.A(n708),
	.B1(FE_OFN62_n4016),
	.B2(n38),
	.ZN(n1715));
   NAND2_X1 U1213 (.A1(REGISTERS[608]),
	.A2(FE_OFN62_n4016),
	.ZN(n708));
   OAI21_X1 U1214 (.A(n710),
	.B1(FE_OFN62_n4016),
	.B2(n42),
	.ZN(n1717));
   NAND2_X1 U1215 (.A1(REGISTERS[610]),
	.A2(FE_OFN62_n4016),
	.ZN(n710));
   OAI21_X1 U1216 (.A(n713),
	.B1(n4016),
	.B2(n48),
	.ZN(n1720));
   NAND2_X1 U1217 (.A1(REGISTERS[613]),
	.A2(n4016),
	.ZN(n713));
   OAI21_X1 U1218 (.A(n714),
	.B1(FE_OFN62_n4016),
	.B2(n50),
	.ZN(n1721));
   NAND2_X1 U1219 (.A1(REGISTERS[614]),
	.A2(FE_OFN62_n4016),
	.ZN(n714));
   OAI21_X1 U1220 (.A(n721),
	.B1(FE_OFN62_n4016),
	.B2(n64),
	.ZN(n1728));
   NAND2_X1 U1221 (.A1(REGISTERS[621]),
	.A2(FE_OFN62_n4016),
	.ZN(n721));
   OAI21_X1 U1222 (.A(n724),
	.B1(n4016),
	.B2(n70),
	.ZN(n1731));
   NAND2_X1 U1223 (.A1(REGISTERS[624]),
	.A2(n4016),
	.ZN(n724));
   OAI21_X1 U1224 (.A(n725),
	.B1(FE_OFN62_n4016),
	.B2(n72),
	.ZN(n1732));
   NAND2_X1 U1225 (.A1(REGISTERS[625]),
	.A2(FE_OFN62_n4016),
	.ZN(n725));
   OAI21_X1 U1226 (.A(n726),
	.B1(FE_OFN62_n4016),
	.B2(n74),
	.ZN(n1733));
   NAND2_X1 U1227 (.A1(REGISTERS[626]),
	.A2(FE_OFN62_n4016),
	.ZN(n726));
   OAI21_X1 U1228 (.A(n727),
	.B1(FE_OFN62_n4016),
	.B2(n76),
	.ZN(n1734));
   NAND2_X1 U1229 (.A1(REGISTERS[627]),
	.A2(FE_OFN62_n4016),
	.ZN(n727));
   OAI21_X1 U1230 (.A(n728),
	.B1(FE_OFN62_n4016),
	.B2(n78),
	.ZN(n1735));
   NAND2_X1 U1231 (.A1(REGISTERS[628]),
	.A2(FE_OFN62_n4016),
	.ZN(n728));
   OAI21_X1 U1232 (.A(n729),
	.B1(FE_OFN62_n4016),
	.B2(n80),
	.ZN(n1736));
   NAND2_X1 U1233 (.A1(REGISTERS[629]),
	.A2(FE_OFN62_n4016),
	.ZN(n729));
   OAI21_X1 U1234 (.A(n730),
	.B1(FE_OFN62_n4016),
	.B2(n82),
	.ZN(n1737));
   NAND2_X1 U1235 (.A1(REGISTERS[630]),
	.A2(FE_OFN62_n4016),
	.ZN(n730));
   OAI21_X1 U1236 (.A(n731),
	.B1(FE_OFN62_n4016),
	.B2(n84),
	.ZN(n1738));
   NAND2_X1 U1237 (.A1(REGISTERS[631]),
	.A2(FE_OFN62_n4016),
	.ZN(n731));
   OAI21_X1 U1238 (.A(n732),
	.B1(FE_OFN62_n4016),
	.B2(n86),
	.ZN(n1739));
   NAND2_X1 U1239 (.A1(REGISTERS[632]),
	.A2(FE_OFN62_n4016),
	.ZN(n732));
   OAI21_X1 U1240 (.A(n733),
	.B1(FE_OFN62_n4016),
	.B2(n88),
	.ZN(n1740));
   NAND2_X1 U1241 (.A1(REGISTERS[633]),
	.A2(FE_OFN62_n4016),
	.ZN(n733));
   OAI21_X1 U1242 (.A(n734),
	.B1(FE_OFN62_n4016),
	.B2(n90),
	.ZN(n1741));
   NAND2_X1 U1243 (.A1(REGISTERS[634]),
	.A2(FE_OFN62_n4016),
	.ZN(n734));
   OAI21_X1 U1244 (.A(n735),
	.B1(FE_OFN62_n4016),
	.B2(n92),
	.ZN(n1742));
   NAND2_X1 U1245 (.A1(REGISTERS[635]),
	.A2(FE_OFN62_n4016),
	.ZN(n735));
   OAI21_X1 U1246 (.A(n736),
	.B1(FE_OFN62_n4016),
	.B2(n94),
	.ZN(n1743));
   NAND2_X1 U1247 (.A1(REGISTERS[636]),
	.A2(FE_OFN62_n4016),
	.ZN(n736));
   OAI21_X1 U1248 (.A(n741),
	.B1(n4015),
	.B2(n38),
	.ZN(n1747));
   NAND2_X1 U1249 (.A1(REGISTERS[640]),
	.A2(n4015),
	.ZN(n741));
   OAI21_X1 U1250 (.A(n743),
	.B1(FE_OFN74_n4015),
	.B2(n42),
	.ZN(n1749));
   NAND2_X1 U1251 (.A1(REGISTERS[642]),
	.A2(FE_OFN74_n4015),
	.ZN(n743));
   OAI21_X1 U1252 (.A(n746),
	.B1(FE_OFN74_n4015),
	.B2(n48),
	.ZN(n1752));
   NAND2_X1 U1253 (.A1(REGISTERS[645]),
	.A2(FE_OFN74_n4015),
	.ZN(n746));
   OAI21_X1 U1254 (.A(n747),
	.B1(n4015),
	.B2(n50),
	.ZN(n1753));
   NAND2_X1 U1255 (.A1(REGISTERS[646]),
	.A2(n4015),
	.ZN(n747));
   OAI21_X1 U1256 (.A(n754),
	.B1(n4015),
	.B2(n64),
	.ZN(n1760));
   NAND2_X1 U1257 (.A1(REGISTERS[653]),
	.A2(n4015),
	.ZN(n754));
   OAI21_X1 U1258 (.A(n757),
	.B1(FE_OFN74_n4015),
	.B2(n70),
	.ZN(n1763));
   NAND2_X1 U1259 (.A1(REGISTERS[656]),
	.A2(FE_OFN74_n4015),
	.ZN(n757));
   OAI21_X1 U1260 (.A(n758),
	.B1(FE_OFN74_n4015),
	.B2(n72),
	.ZN(n1764));
   NAND2_X1 U1261 (.A1(REGISTERS[657]),
	.A2(FE_OFN74_n4015),
	.ZN(n758));
   OAI21_X1 U1262 (.A(n759),
	.B1(n4015),
	.B2(n74),
	.ZN(n1765));
   NAND2_X1 U1263 (.A1(REGISTERS[658]),
	.A2(n4015),
	.ZN(n759));
   OAI21_X1 U1264 (.A(n760),
	.B1(FE_OFN74_n4015),
	.B2(n76),
	.ZN(n1766));
   NAND2_X1 U1265 (.A1(REGISTERS[659]),
	.A2(FE_OFN74_n4015),
	.ZN(n760));
   OAI21_X1 U1266 (.A(n761),
	.B1(n4015),
	.B2(n78),
	.ZN(n1767));
   NAND2_X1 U1267 (.A1(REGISTERS[660]),
	.A2(n4015),
	.ZN(n761));
   OAI21_X1 U1268 (.A(n762),
	.B1(FE_OFN74_n4015),
	.B2(n80),
	.ZN(n1768));
   NAND2_X1 U1269 (.A1(REGISTERS[661]),
	.A2(FE_OFN74_n4015),
	.ZN(n762));
   OAI21_X1 U1270 (.A(n763),
	.B1(FE_OFN74_n4015),
	.B2(n82),
	.ZN(n1769));
   NAND2_X1 U1271 (.A1(REGISTERS[662]),
	.A2(FE_OFN74_n4015),
	.ZN(n763));
   OAI21_X1 U1272 (.A(n764),
	.B1(FE_OFN74_n4015),
	.B2(n84),
	.ZN(n1770));
   NAND2_X1 U1273 (.A1(REGISTERS[663]),
	.A2(FE_OFN74_n4015),
	.ZN(n764));
   OAI21_X1 U1274 (.A(n765),
	.B1(n4015),
	.B2(n86),
	.ZN(n1771));
   NAND2_X1 U1275 (.A1(REGISTERS[664]),
	.A2(n4015),
	.ZN(n765));
   OAI21_X1 U1276 (.A(n766),
	.B1(FE_OFN74_n4015),
	.B2(n88),
	.ZN(n1772));
   NAND2_X1 U1277 (.A1(REGISTERS[665]),
	.A2(FE_OFN74_n4015),
	.ZN(n766));
   OAI21_X1 U1278 (.A(n767),
	.B1(n4015),
	.B2(n90),
	.ZN(n1773));
   NAND2_X1 U1279 (.A1(REGISTERS[666]),
	.A2(n4015),
	.ZN(n767));
   OAI21_X1 U1280 (.A(n768),
	.B1(FE_OFN74_n4015),
	.B2(n92),
	.ZN(n1774));
   NAND2_X1 U1281 (.A1(REGISTERS[667]),
	.A2(FE_OFN74_n4015),
	.ZN(n768));
   OAI21_X1 U1282 (.A(n769),
	.B1(FE_OFN74_n4015),
	.B2(n94),
	.ZN(n1775));
   NAND2_X1 U1283 (.A1(REGISTERS[668]),
	.A2(FE_OFN74_n4015),
	.ZN(n769));
   OAI21_X1 U1284 (.A(n774),
	.B1(n4014),
	.B2(n38),
	.ZN(n1779));
   NAND2_X1 U1285 (.A1(REGISTERS[672]),
	.A2(n4014),
	.ZN(n774));
   OAI21_X1 U1286 (.A(n776),
	.B1(FE_OFN78_n4014),
	.B2(n42),
	.ZN(n1781));
   NAND2_X1 U1287 (.A1(REGISTERS[674]),
	.A2(FE_OFN78_n4014),
	.ZN(n776));
   OAI21_X1 U1288 (.A(n779),
	.B1(FE_OFN78_n4014),
	.B2(n48),
	.ZN(n1784));
   NAND2_X1 U1289 (.A1(REGISTERS[677]),
	.A2(FE_OFN78_n4014),
	.ZN(n779));
   OAI21_X1 U1290 (.A(n780),
	.B1(n4014),
	.B2(n50),
	.ZN(n1785));
   NAND2_X1 U1291 (.A1(REGISTERS[678]),
	.A2(n4014),
	.ZN(n780));
   OAI21_X1 U1292 (.A(n787),
	.B1(n4014),
	.B2(n64),
	.ZN(n1792));
   NAND2_X1 U1293 (.A1(REGISTERS[685]),
	.A2(n4014),
	.ZN(n787));
   OAI21_X1 U1294 (.A(n790),
	.B1(FE_OFN78_n4014),
	.B2(n70),
	.ZN(n1795));
   NAND2_X1 U1295 (.A1(REGISTERS[688]),
	.A2(FE_OFN78_n4014),
	.ZN(n790));
   OAI21_X1 U1296 (.A(n791),
	.B1(FE_OFN78_n4014),
	.B2(n72),
	.ZN(n1796));
   NAND2_X1 U1297 (.A1(REGISTERS[689]),
	.A2(FE_OFN78_n4014),
	.ZN(n791));
   OAI21_X1 U1298 (.A(n792),
	.B1(n4014),
	.B2(n74),
	.ZN(n1797));
   NAND2_X1 U1299 (.A1(REGISTERS[690]),
	.A2(n4014),
	.ZN(n792));
   OAI21_X1 U1300 (.A(n793),
	.B1(FE_OFN78_n4014),
	.B2(n76),
	.ZN(n1798));
   NAND2_X1 U1301 (.A1(REGISTERS[691]),
	.A2(FE_OFN78_n4014),
	.ZN(n793));
   OAI21_X1 U1302 (.A(n794),
	.B1(FE_OFN78_n4014),
	.B2(n78),
	.ZN(n1799));
   NAND2_X1 U1303 (.A1(REGISTERS[692]),
	.A2(FE_OFN78_n4014),
	.ZN(n794));
   OAI21_X1 U1304 (.A(n795),
	.B1(FE_OFN78_n4014),
	.B2(n80),
	.ZN(n1800));
   NAND2_X1 U1305 (.A1(REGISTERS[693]),
	.A2(FE_OFN78_n4014),
	.ZN(n795));
   OAI21_X1 U1306 (.A(n796),
	.B1(FE_OFN78_n4014),
	.B2(n82),
	.ZN(n1801));
   NAND2_X1 U1307 (.A1(REGISTERS[694]),
	.A2(FE_OFN78_n4014),
	.ZN(n796));
   OAI21_X1 U1308 (.A(n797),
	.B1(FE_OFN78_n4014),
	.B2(n84),
	.ZN(n1802));
   NAND2_X1 U1309 (.A1(REGISTERS[695]),
	.A2(FE_OFN78_n4014),
	.ZN(n797));
   OAI21_X1 U1310 (.A(n798),
	.B1(FE_OFN78_n4014),
	.B2(n86),
	.ZN(n1803));
   NAND2_X1 U1311 (.A1(REGISTERS[696]),
	.A2(FE_OFN78_n4014),
	.ZN(n798));
   OAI21_X1 U1312 (.A(n799),
	.B1(FE_OFN78_n4014),
	.B2(n88),
	.ZN(n1804));
   NAND2_X1 U1313 (.A1(REGISTERS[697]),
	.A2(FE_OFN78_n4014),
	.ZN(n799));
   OAI21_X1 U1314 (.A(n800),
	.B1(FE_OFN78_n4014),
	.B2(n90),
	.ZN(n1805));
   NAND2_X1 U1315 (.A1(REGISTERS[698]),
	.A2(FE_OFN78_n4014),
	.ZN(n800));
   OAI21_X1 U1316 (.A(n801),
	.B1(FE_OFN78_n4014),
	.B2(n92),
	.ZN(n1806));
   NAND2_X1 U1317 (.A1(REGISTERS[699]),
	.A2(FE_OFN78_n4014),
	.ZN(n801));
   OAI21_X1 U1318 (.A(n802),
	.B1(FE_OFN78_n4014),
	.B2(n94),
	.ZN(n1807));
   NAND2_X1 U1319 (.A1(REGISTERS[700]),
	.A2(FE_OFN78_n4014),
	.ZN(n802));
   OAI21_X1 U1320 (.A(n807),
	.B1(n4013),
	.B2(n38),
	.ZN(n1811));
   NAND2_X1 U1321 (.A1(REGISTERS[704]),
	.A2(n4013),
	.ZN(n807));
   OAI21_X1 U1322 (.A(n809),
	.B1(FE_OFN76_n4013),
	.B2(n42),
	.ZN(n1813));
   NAND2_X1 U1323 (.A1(REGISTERS[706]),
	.A2(FE_OFN76_n4013),
	.ZN(n809));
   OAI21_X1 U1324 (.A(n812),
	.B1(FE_OFN76_n4013),
	.B2(n48),
	.ZN(n1816));
   NAND2_X1 U1325 (.A1(REGISTERS[709]),
	.A2(FE_OFN76_n4013),
	.ZN(n812));
   OAI21_X1 U1326 (.A(n813),
	.B1(n4013),
	.B2(n50),
	.ZN(n1817));
   NAND2_X1 U1327 (.A1(REGISTERS[710]),
	.A2(n4013),
	.ZN(n813));
   OAI21_X1 U1328 (.A(n820),
	.B1(n4013),
	.B2(n64),
	.ZN(n1824));
   NAND2_X1 U1329 (.A1(REGISTERS[717]),
	.A2(n4013),
	.ZN(n820));
   OAI21_X1 U1330 (.A(n823),
	.B1(FE_OFN76_n4013),
	.B2(n70),
	.ZN(n1827));
   NAND2_X1 U1331 (.A1(REGISTERS[720]),
	.A2(FE_OFN76_n4013),
	.ZN(n823));
   OAI21_X1 U1332 (.A(n824),
	.B1(FE_OFN76_n4013),
	.B2(n72),
	.ZN(n1828));
   NAND2_X1 U1333 (.A1(REGISTERS[721]),
	.A2(FE_OFN76_n4013),
	.ZN(n824));
   OAI21_X1 U1334 (.A(n825),
	.B1(n4013),
	.B2(n74),
	.ZN(n1829));
   NAND2_X1 U1335 (.A1(REGISTERS[722]),
	.A2(n4013),
	.ZN(n825));
   OAI21_X1 U1336 (.A(n826),
	.B1(FE_OFN76_n4013),
	.B2(n76),
	.ZN(n1830));
   NAND2_X1 U1337 (.A1(REGISTERS[723]),
	.A2(FE_OFN76_n4013),
	.ZN(n826));
   OAI21_X1 U1338 (.A(n827),
	.B1(n4013),
	.B2(n78),
	.ZN(n1831));
   NAND2_X1 U1339 (.A1(REGISTERS[724]),
	.A2(n4013),
	.ZN(n827));
   OAI21_X1 U1340 (.A(n828),
	.B1(FE_OFN76_n4013),
	.B2(n80),
	.ZN(n1832));
   NAND2_X1 U1341 (.A1(REGISTERS[725]),
	.A2(FE_OFN76_n4013),
	.ZN(n828));
   OAI21_X1 U1342 (.A(n829),
	.B1(FE_OFN76_n4013),
	.B2(n82),
	.ZN(n1833));
   NAND2_X1 U1343 (.A1(REGISTERS[726]),
	.A2(FE_OFN76_n4013),
	.ZN(n829));
   OAI21_X1 U1344 (.A(n830),
	.B1(FE_OFN76_n4013),
	.B2(n84),
	.ZN(n1834));
   NAND2_X1 U1345 (.A1(REGISTERS[727]),
	.A2(FE_OFN76_n4013),
	.ZN(n830));
   OAI21_X1 U1346 (.A(n831),
	.B1(n4013),
	.B2(n86),
	.ZN(n1835));
   NAND2_X1 U1347 (.A1(REGISTERS[728]),
	.A2(n4013),
	.ZN(n831));
   OAI21_X1 U1348 (.A(n832),
	.B1(FE_OFN76_n4013),
	.B2(n88),
	.ZN(n1836));
   NAND2_X1 U1349 (.A1(REGISTERS[729]),
	.A2(FE_OFN76_n4013),
	.ZN(n832));
   OAI21_X1 U1350 (.A(n833),
	.B1(n4013),
	.B2(n90),
	.ZN(n1837));
   NAND2_X1 U1351 (.A1(REGISTERS[730]),
	.A2(n4013),
	.ZN(n833));
   OAI21_X1 U1352 (.A(n834),
	.B1(FE_OFN76_n4013),
	.B2(n92),
	.ZN(n1838));
   NAND2_X1 U1353 (.A1(REGISTERS[731]),
	.A2(FE_OFN76_n4013),
	.ZN(n834));
   OAI21_X1 U1354 (.A(n835),
	.B1(FE_OFN76_n4013),
	.B2(n94),
	.ZN(n1839));
   NAND2_X1 U1355 (.A1(REGISTERS[732]),
	.A2(FE_OFN76_n4013),
	.ZN(n835));
   OAI21_X1 U1356 (.A(n840),
	.B1(n4012),
	.B2(n38),
	.ZN(n1843));
   NAND2_X1 U1357 (.A1(REGISTERS[736]),
	.A2(n4012),
	.ZN(n840));
   OAI21_X1 U1358 (.A(n842),
	.B1(FE_OFN64_n4012),
	.B2(n42),
	.ZN(n1845));
   NAND2_X1 U1359 (.A1(REGISTERS[738]),
	.A2(FE_OFN64_n4012),
	.ZN(n842));
   OAI21_X1 U1360 (.A(n845),
	.B1(FE_OFN64_n4012),
	.B2(n48),
	.ZN(n1848));
   NAND2_X1 U1361 (.A1(REGISTERS[741]),
	.A2(FE_OFN64_n4012),
	.ZN(n845));
   OAI21_X1 U1362 (.A(n846),
	.B1(n4012),
	.B2(n50),
	.ZN(n1849));
   NAND2_X1 U1363 (.A1(REGISTERS[742]),
	.A2(n4012),
	.ZN(n846));
   OAI21_X1 U1364 (.A(n853),
	.B1(n4012),
	.B2(n64),
	.ZN(n1856));
   NAND2_X1 U1365 (.A1(REGISTERS[749]),
	.A2(n4012),
	.ZN(n853));
   OAI21_X1 U1366 (.A(n856),
	.B1(FE_OFN64_n4012),
	.B2(n70),
	.ZN(n1859));
   NAND2_X1 U1367 (.A1(REGISTERS[752]),
	.A2(FE_OFN64_n4012),
	.ZN(n856));
   OAI21_X1 U1368 (.A(n857),
	.B1(FE_OFN64_n4012),
	.B2(n72),
	.ZN(n1860));
   NAND2_X1 U1369 (.A1(REGISTERS[753]),
	.A2(FE_OFN64_n4012),
	.ZN(n857));
   OAI21_X1 U1370 (.A(n858),
	.B1(n4012),
	.B2(n74),
	.ZN(n1861));
   NAND2_X1 U1371 (.A1(REGISTERS[754]),
	.A2(n4012),
	.ZN(n858));
   OAI21_X1 U1372 (.A(n859),
	.B1(FE_OFN64_n4012),
	.B2(n76),
	.ZN(n1862));
   NAND2_X1 U1373 (.A1(REGISTERS[755]),
	.A2(FE_OFN64_n4012),
	.ZN(n859));
   OAI21_X1 U1374 (.A(n860),
	.B1(FE_OFN64_n4012),
	.B2(n78),
	.ZN(n1863));
   NAND2_X1 U1375 (.A1(REGISTERS[756]),
	.A2(FE_OFN64_n4012),
	.ZN(n860));
   OAI21_X1 U1376 (.A(n861),
	.B1(FE_OFN64_n4012),
	.B2(n80),
	.ZN(n1864));
   NAND2_X1 U1377 (.A1(REGISTERS[757]),
	.A2(FE_OFN64_n4012),
	.ZN(n861));
   OAI21_X1 U1378 (.A(n862),
	.B1(FE_OFN64_n4012),
	.B2(n82),
	.ZN(n1865));
   NAND2_X1 U1379 (.A1(REGISTERS[758]),
	.A2(FE_OFN64_n4012),
	.ZN(n862));
   OAI21_X1 U1380 (.A(n863),
	.B1(FE_OFN64_n4012),
	.B2(n84),
	.ZN(n1866));
   NAND2_X1 U1381 (.A1(REGISTERS[759]),
	.A2(FE_OFN64_n4012),
	.ZN(n863));
   OAI21_X1 U1382 (.A(n864),
	.B1(FE_OFN64_n4012),
	.B2(n86),
	.ZN(n1867));
   NAND2_X1 U1383 (.A1(REGISTERS[760]),
	.A2(FE_OFN64_n4012),
	.ZN(n864));
   OAI21_X1 U1384 (.A(n865),
	.B1(FE_OFN64_n4012),
	.B2(n88),
	.ZN(n1868));
   NAND2_X1 U1385 (.A1(REGISTERS[761]),
	.A2(FE_OFN64_n4012),
	.ZN(n865));
   OAI21_X1 U1386 (.A(n866),
	.B1(FE_OFN64_n4012),
	.B2(n90),
	.ZN(n1869));
   NAND2_X1 U1387 (.A1(REGISTERS[762]),
	.A2(FE_OFN64_n4012),
	.ZN(n866));
   OAI21_X1 U1388 (.A(n867),
	.B1(FE_OFN64_n4012),
	.B2(n92),
	.ZN(n1870));
   NAND2_X1 U1389 (.A1(REGISTERS[763]),
	.A2(FE_OFN64_n4012),
	.ZN(n867));
   OAI21_X1 U1390 (.A(n868),
	.B1(FE_OFN64_n4012),
	.B2(n94),
	.ZN(n1871));
   NAND2_X1 U1391 (.A1(REGISTERS[764]),
	.A2(FE_OFN64_n4012),
	.ZN(n868));
   OAI21_X1 U1392 (.A(n873),
	.B1(n4011),
	.B2(n38),
	.ZN(n1875));
   NAND2_X1 U1393 (.A1(REGISTERS[768]),
	.A2(n4011),
	.ZN(n873));
   OAI21_X1 U1394 (.A(n875),
	.B1(FE_OFN68_n4011),
	.B2(n42),
	.ZN(n1877));
   NAND2_X1 U1395 (.A1(REGISTERS[770]),
	.A2(FE_OFN68_n4011),
	.ZN(n875));
   OAI21_X1 U1396 (.A(n878),
	.B1(FE_OFN68_n4011),
	.B2(n48),
	.ZN(n1880));
   NAND2_X1 U1397 (.A1(REGISTERS[773]),
	.A2(FE_OFN68_n4011),
	.ZN(n878));
   OAI21_X1 U1398 (.A(n879),
	.B1(n4011),
	.B2(n50),
	.ZN(n1881));
   NAND2_X1 U1399 (.A1(REGISTERS[774]),
	.A2(n4011),
	.ZN(n879));
   OAI21_X1 U1400 (.A(n880),
	.B1(FE_OFN68_n4011),
	.B2(n52),
	.ZN(n1882));
   NAND2_X1 U1401 (.A1(REGISTERS[775]),
	.A2(FE_OFN68_n4011),
	.ZN(n880));
   OAI21_X1 U1402 (.A(n881),
	.B1(n4011),
	.B2(n54),
	.ZN(n1883));
   NAND2_X1 U1403 (.A1(REGISTERS[776]),
	.A2(n4011),
	.ZN(n881));
   OAI21_X1 U1404 (.A(n882),
	.B1(FE_OFN68_n4011),
	.B2(n56),
	.ZN(n1884));
   NAND2_X1 U1405 (.A1(REGISTERS[777]),
	.A2(FE_OFN68_n4011),
	.ZN(n882));
   OAI21_X1 U1406 (.A(n883),
	.B1(n4011),
	.B2(n58),
	.ZN(n1885));
   NAND2_X1 U1407 (.A1(REGISTERS[778]),
	.A2(n4011),
	.ZN(n883));
   OAI21_X1 U1408 (.A(n884),
	.B1(FE_OFN68_n4011),
	.B2(n60),
	.ZN(n1886));
   NAND2_X1 U1409 (.A1(REGISTERS[779]),
	.A2(FE_OFN68_n4011),
	.ZN(n884));
   OAI21_X1 U1410 (.A(n885),
	.B1(n4011),
	.B2(n62),
	.ZN(n1887));
   NAND2_X1 U1411 (.A1(REGISTERS[780]),
	.A2(n4011),
	.ZN(n885));
   OAI21_X1 U1412 (.A(n886),
	.B1(n4011),
	.B2(n64),
	.ZN(n1888));
   NAND2_X1 U1413 (.A1(REGISTERS[781]),
	.A2(n4011),
	.ZN(n886));
   OAI21_X1 U1414 (.A(n887),
	.B1(FE_OFN68_n4011),
	.B2(n66),
	.ZN(n1889));
   NAND2_X1 U1415 (.A1(REGISTERS[782]),
	.A2(FE_OFN68_n4011),
	.ZN(n887));
   OAI21_X1 U1416 (.A(n888),
	.B1(FE_OFN68_n4011),
	.B2(n68),
	.ZN(n1890));
   NAND2_X1 U1417 (.A1(REGISTERS[783]),
	.A2(FE_OFN68_n4011),
	.ZN(n888));
   OAI21_X1 U1418 (.A(n889),
	.B1(FE_OFN68_n4011),
	.B2(n70),
	.ZN(n1891));
   NAND2_X1 U1419 (.A1(REGISTERS[784]),
	.A2(FE_OFN68_n4011),
	.ZN(n889));
   OAI21_X1 U1420 (.A(n890),
	.B1(FE_OFN68_n4011),
	.B2(n72),
	.ZN(n1892));
   NAND2_X1 U1421 (.A1(REGISTERS[785]),
	.A2(FE_OFN68_n4011),
	.ZN(n890));
   OAI21_X1 U1422 (.A(n891),
	.B1(n4011),
	.B2(n74),
	.ZN(n1893));
   NAND2_X1 U1423 (.A1(REGISTERS[786]),
	.A2(n4011),
	.ZN(n891));
   OAI21_X1 U1424 (.A(n892),
	.B1(FE_OFN68_n4011),
	.B2(n76),
	.ZN(n1894));
   NAND2_X1 U1425 (.A1(REGISTERS[787]),
	.A2(FE_OFN68_n4011),
	.ZN(n892));
   OAI21_X1 U1426 (.A(n893),
	.B1(n4011),
	.B2(n78),
	.ZN(n1895));
   NAND2_X1 U1427 (.A1(REGISTERS[788]),
	.A2(n4011),
	.ZN(n893));
   OAI21_X1 U1428 (.A(n894),
	.B1(FE_OFN68_n4011),
	.B2(n80),
	.ZN(n1896));
   NAND2_X1 U1429 (.A1(REGISTERS[789]),
	.A2(FE_OFN68_n4011),
	.ZN(n894));
   OAI21_X1 U1430 (.A(n895),
	.B1(FE_OFN68_n4011),
	.B2(n82),
	.ZN(n1897));
   NAND2_X1 U1431 (.A1(REGISTERS[790]),
	.A2(FE_OFN68_n4011),
	.ZN(n895));
   OAI21_X1 U1432 (.A(n896),
	.B1(FE_OFN68_n4011),
	.B2(n84),
	.ZN(n1898));
   NAND2_X1 U1433 (.A1(REGISTERS[791]),
	.A2(FE_OFN68_n4011),
	.ZN(n896));
   OAI21_X1 U1434 (.A(n897),
	.B1(n4011),
	.B2(n86),
	.ZN(n1899));
   NAND2_X1 U1435 (.A1(REGISTERS[792]),
	.A2(n4011),
	.ZN(n897));
   OAI21_X1 U1436 (.A(n898),
	.B1(FE_OFN68_n4011),
	.B2(n88),
	.ZN(n1900));
   NAND2_X1 U1437 (.A1(REGISTERS[793]),
	.A2(FE_OFN68_n4011),
	.ZN(n898));
   OAI21_X1 U1438 (.A(n899),
	.B1(n4011),
	.B2(n90),
	.ZN(n1901));
   NAND2_X1 U1439 (.A1(REGISTERS[794]),
	.A2(n4011),
	.ZN(n899));
   OAI21_X1 U1440 (.A(n900),
	.B1(FE_OFN68_n4011),
	.B2(n92),
	.ZN(n1902));
   NAND2_X1 U1441 (.A1(REGISTERS[795]),
	.A2(FE_OFN68_n4011),
	.ZN(n900));
   OAI21_X1 U1442 (.A(n901),
	.B1(FE_OFN68_n4011),
	.B2(n94),
	.ZN(n1903));
   NAND2_X1 U1443 (.A1(REGISTERS[796]),
	.A2(FE_OFN68_n4011),
	.ZN(n901));
   OAI21_X1 U1444 (.A(n907),
	.B1(n4010),
	.B2(n38),
	.ZN(n1907));
   NAND2_X1 U1445 (.A1(REGISTERS[800]),
	.A2(n4010),
	.ZN(n907));
   OAI21_X1 U1446 (.A(n909),
	.B1(FE_OFN88_n4010),
	.B2(n42),
	.ZN(n1909));
   NAND2_X1 U1447 (.A1(REGISTERS[802]),
	.A2(FE_OFN88_n4010),
	.ZN(n909));
   OAI21_X1 U1448 (.A(n912),
	.B1(FE_OFN88_n4010),
	.B2(n48),
	.ZN(n1912));
   NAND2_X1 U1449 (.A1(REGISTERS[805]),
	.A2(FE_OFN88_n4010),
	.ZN(n912));
   OAI21_X1 U1450 (.A(n913),
	.B1(n4010),
	.B2(n50),
	.ZN(n1913));
   NAND2_X1 U1451 (.A1(REGISTERS[806]),
	.A2(n4010),
	.ZN(n913));
   OAI21_X1 U1452 (.A(n914),
	.B1(FE_OFN88_n4010),
	.B2(n52),
	.ZN(n1914));
   NAND2_X1 U1453 (.A1(REGISTERS[807]),
	.A2(FE_OFN88_n4010),
	.ZN(n914));
   OAI21_X1 U1454 (.A(n915),
	.B1(n4010),
	.B2(n54),
	.ZN(n1915));
   NAND2_X1 U1455 (.A1(REGISTERS[808]),
	.A2(n4010),
	.ZN(n915));
   OAI21_X1 U1456 (.A(n916),
	.B1(FE_OFN88_n4010),
	.B2(n56),
	.ZN(n1916));
   NAND2_X1 U1457 (.A1(REGISTERS[809]),
	.A2(FE_OFN88_n4010),
	.ZN(n916));
   OAI21_X1 U1458 (.A(n917),
	.B1(n4010),
	.B2(n58),
	.ZN(n1917));
   NAND2_X1 U1459 (.A1(REGISTERS[810]),
	.A2(n4010),
	.ZN(n917));
   OAI21_X1 U1460 (.A(n918),
	.B1(FE_OFN88_n4010),
	.B2(n60),
	.ZN(n1918));
   NAND2_X1 U1461 (.A1(REGISTERS[811]),
	.A2(FE_OFN88_n4010),
	.ZN(n918));
   OAI21_X1 U1462 (.A(n919),
	.B1(n4010),
	.B2(n62),
	.ZN(n1919));
   NAND2_X1 U1463 (.A1(REGISTERS[812]),
	.A2(n4010),
	.ZN(n919));
   OAI21_X1 U1464 (.A(n920),
	.B1(n4010),
	.B2(n64),
	.ZN(n1920));
   NAND2_X1 U1465 (.A1(REGISTERS[813]),
	.A2(n4010),
	.ZN(n920));
   OAI21_X1 U1466 (.A(n921),
	.B1(FE_OFN88_n4010),
	.B2(n66),
	.ZN(n1921));
   NAND2_X1 U1467 (.A1(REGISTERS[814]),
	.A2(FE_OFN88_n4010),
	.ZN(n921));
   OAI21_X1 U1468 (.A(n922),
	.B1(FE_OFN88_n4010),
	.B2(n68),
	.ZN(n1922));
   NAND2_X1 U1469 (.A1(REGISTERS[815]),
	.A2(FE_OFN88_n4010),
	.ZN(n922));
   OAI21_X1 U1470 (.A(n923),
	.B1(FE_OFN88_n4010),
	.B2(n70),
	.ZN(n1923));
   NAND2_X1 U1471 (.A1(REGISTERS[816]),
	.A2(FE_OFN88_n4010),
	.ZN(n923));
   OAI21_X1 U1472 (.A(n924),
	.B1(FE_OFN88_n4010),
	.B2(n72),
	.ZN(n1924));
   NAND2_X1 U1473 (.A1(REGISTERS[817]),
	.A2(FE_OFN88_n4010),
	.ZN(n924));
   OAI21_X1 U1474 (.A(n925),
	.B1(n4010),
	.B2(n74),
	.ZN(n1925));
   NAND2_X1 U1475 (.A1(REGISTERS[818]),
	.A2(n4010),
	.ZN(n925));
   OAI21_X1 U1476 (.A(n926),
	.B1(FE_OFN88_n4010),
	.B2(n76),
	.ZN(n1926));
   NAND2_X1 U1477 (.A1(REGISTERS[819]),
	.A2(FE_OFN88_n4010),
	.ZN(n926));
   OAI21_X1 U1478 (.A(n927),
	.B1(n4010),
	.B2(n78),
	.ZN(n1927));
   NAND2_X1 U1479 (.A1(REGISTERS[820]),
	.A2(n4010),
	.ZN(n927));
   OAI21_X1 U1480 (.A(n928),
	.B1(FE_OFN88_n4010),
	.B2(n80),
	.ZN(n1928));
   NAND2_X1 U1481 (.A1(REGISTERS[821]),
	.A2(FE_OFN88_n4010),
	.ZN(n928));
   OAI21_X1 U1482 (.A(n929),
	.B1(FE_OFN88_n4010),
	.B2(n82),
	.ZN(n1929));
   NAND2_X1 U1483 (.A1(REGISTERS[822]),
	.A2(FE_OFN88_n4010),
	.ZN(n929));
   OAI21_X1 U1484 (.A(n930),
	.B1(FE_OFN88_n4010),
	.B2(n84),
	.ZN(n1930));
   NAND2_X1 U1485 (.A1(REGISTERS[823]),
	.A2(FE_OFN88_n4010),
	.ZN(n930));
   OAI21_X1 U1486 (.A(n931),
	.B1(n4010),
	.B2(n86),
	.ZN(n1931));
   NAND2_X1 U1487 (.A1(REGISTERS[824]),
	.A2(n4010),
	.ZN(n931));
   OAI21_X1 U1488 (.A(n932),
	.B1(FE_OFN88_n4010),
	.B2(n88),
	.ZN(n1932));
   NAND2_X1 U1489 (.A1(REGISTERS[825]),
	.A2(FE_OFN88_n4010),
	.ZN(n932));
   OAI21_X1 U1490 (.A(n933),
	.B1(n4010),
	.B2(n90),
	.ZN(n1933));
   NAND2_X1 U1491 (.A1(REGISTERS[826]),
	.A2(n4010),
	.ZN(n933));
   OAI21_X1 U1492 (.A(n934),
	.B1(FE_OFN88_n4010),
	.B2(n92),
	.ZN(n1934));
   NAND2_X1 U1493 (.A1(REGISTERS[827]),
	.A2(FE_OFN88_n4010),
	.ZN(n934));
   OAI21_X1 U1494 (.A(n935),
	.B1(FE_OFN88_n4010),
	.B2(n94),
	.ZN(n1935));
   NAND2_X1 U1495 (.A1(REGISTERS[828]),
	.A2(FE_OFN88_n4010),
	.ZN(n935));
   OAI21_X1 U1496 (.A(n940),
	.B1(n4009),
	.B2(n38),
	.ZN(n1939));
   NAND2_X1 U1497 (.A1(REGISTERS[832]),
	.A2(n4009),
	.ZN(n940));
   OAI21_X1 U1498 (.A(n942),
	.B1(FE_OFN73_n4009),
	.B2(n42),
	.ZN(n1941));
   NAND2_X1 U1499 (.A1(REGISTERS[834]),
	.A2(FE_OFN73_n4009),
	.ZN(n942));
   OAI21_X1 U1500 (.A(n945),
	.B1(FE_OFN73_n4009),
	.B2(n48),
	.ZN(n1944));
   NAND2_X1 U1501 (.A1(REGISTERS[837]),
	.A2(FE_OFN73_n4009),
	.ZN(n945));
   OAI21_X1 U1502 (.A(n946),
	.B1(n4009),
	.B2(n50),
	.ZN(n1945));
   NAND2_X1 U1503 (.A1(REGISTERS[838]),
	.A2(n4009),
	.ZN(n946));
   OAI21_X1 U1504 (.A(n947),
	.B1(FE_OFN73_n4009),
	.B2(n52),
	.ZN(n1946));
   NAND2_X1 U1505 (.A1(REGISTERS[839]),
	.A2(FE_OFN73_n4009),
	.ZN(n947));
   OAI21_X1 U1506 (.A(n948),
	.B1(n4009),
	.B2(n54),
	.ZN(n1947));
   NAND2_X1 U1507 (.A1(REGISTERS[840]),
	.A2(n4009),
	.ZN(n948));
   OAI21_X1 U1508 (.A(n949),
	.B1(FE_OFN73_n4009),
	.B2(n56),
	.ZN(n1948));
   NAND2_X1 U1509 (.A1(REGISTERS[841]),
	.A2(FE_OFN73_n4009),
	.ZN(n949));
   OAI21_X1 U1510 (.A(n950),
	.B1(n4009),
	.B2(n58),
	.ZN(n1949));
   NAND2_X1 U1511 (.A1(REGISTERS[842]),
	.A2(n4009),
	.ZN(n950));
   OAI21_X1 U1512 (.A(n951),
	.B1(FE_OFN73_n4009),
	.B2(n60),
	.ZN(n1950));
   NAND2_X1 U1513 (.A1(REGISTERS[843]),
	.A2(FE_OFN73_n4009),
	.ZN(n951));
   OAI21_X1 U1514 (.A(n952),
	.B1(n4009),
	.B2(n62),
	.ZN(n1951));
   NAND2_X1 U1515 (.A1(REGISTERS[844]),
	.A2(n4009),
	.ZN(n952));
   OAI21_X1 U1516 (.A(n953),
	.B1(n4009),
	.B2(n64),
	.ZN(n1952));
   NAND2_X1 U1517 (.A1(REGISTERS[845]),
	.A2(n4009),
	.ZN(n953));
   OAI21_X1 U1518 (.A(n954),
	.B1(FE_OFN73_n4009),
	.B2(n66),
	.ZN(n1953));
   NAND2_X1 U1519 (.A1(REGISTERS[846]),
	.A2(FE_OFN73_n4009),
	.ZN(n954));
   OAI21_X1 U1520 (.A(n955),
	.B1(FE_OFN73_n4009),
	.B2(n68),
	.ZN(n1954));
   NAND2_X1 U1521 (.A1(REGISTERS[847]),
	.A2(FE_OFN73_n4009),
	.ZN(n955));
   OAI21_X1 U1522 (.A(n956),
	.B1(FE_OFN73_n4009),
	.B2(n70),
	.ZN(n1955));
   NAND2_X1 U1523 (.A1(REGISTERS[848]),
	.A2(FE_OFN73_n4009),
	.ZN(n956));
   OAI21_X1 U1524 (.A(n957),
	.B1(FE_OFN73_n4009),
	.B2(n72),
	.ZN(n1956));
   NAND2_X1 U1525 (.A1(REGISTERS[849]),
	.A2(FE_OFN73_n4009),
	.ZN(n957));
   OAI21_X1 U1526 (.A(n958),
	.B1(n4009),
	.B2(n74),
	.ZN(n1957));
   NAND2_X1 U1527 (.A1(REGISTERS[850]),
	.A2(n4009),
	.ZN(n958));
   OAI21_X1 U1528 (.A(n959),
	.B1(FE_OFN73_n4009),
	.B2(n76),
	.ZN(n1958));
   NAND2_X1 U1529 (.A1(REGISTERS[851]),
	.A2(FE_OFN73_n4009),
	.ZN(n959));
   OAI21_X1 U1530 (.A(n960),
	.B1(n4009),
	.B2(n78),
	.ZN(n1959));
   NAND2_X1 U1531 (.A1(REGISTERS[852]),
	.A2(n4009),
	.ZN(n960));
   OAI21_X1 U1532 (.A(n961),
	.B1(FE_OFN73_n4009),
	.B2(n80),
	.ZN(n1960));
   NAND2_X1 U1533 (.A1(REGISTERS[853]),
	.A2(FE_OFN73_n4009),
	.ZN(n961));
   OAI21_X1 U1534 (.A(n962),
	.B1(FE_OFN73_n4009),
	.B2(n82),
	.ZN(n1961));
   NAND2_X1 U1535 (.A1(REGISTERS[854]),
	.A2(FE_OFN73_n4009),
	.ZN(n962));
   OAI21_X1 U1536 (.A(n963),
	.B1(FE_OFN73_n4009),
	.B2(n84),
	.ZN(n1962));
   NAND2_X1 U1537 (.A1(REGISTERS[855]),
	.A2(FE_OFN73_n4009),
	.ZN(n963));
   OAI21_X1 U1538 (.A(n964),
	.B1(n4009),
	.B2(n86),
	.ZN(n1963));
   NAND2_X1 U1539 (.A1(REGISTERS[856]),
	.A2(n4009),
	.ZN(n964));
   OAI21_X1 U1540 (.A(n965),
	.B1(FE_OFN73_n4009),
	.B2(n88),
	.ZN(n1964));
   NAND2_X1 U1541 (.A1(REGISTERS[857]),
	.A2(FE_OFN73_n4009),
	.ZN(n965));
   OAI21_X1 U1542 (.A(n966),
	.B1(n4009),
	.B2(n90),
	.ZN(n1965));
   NAND2_X1 U1543 (.A1(REGISTERS[858]),
	.A2(n4009),
	.ZN(n966));
   OAI21_X1 U1544 (.A(n967),
	.B1(FE_OFN73_n4009),
	.B2(n92),
	.ZN(n1966));
   NAND2_X1 U1545 (.A1(REGISTERS[859]),
	.A2(FE_OFN73_n4009),
	.ZN(n967));
   OAI21_X1 U1546 (.A(n968),
	.B1(FE_OFN73_n4009),
	.B2(n94),
	.ZN(n1967));
   NAND2_X1 U1547 (.A1(REGISTERS[860]),
	.A2(FE_OFN73_n4009),
	.ZN(n968));
   OAI21_X1 U1548 (.A(n973),
	.B1(n4008),
	.B2(n38),
	.ZN(n1971));
   NAND2_X1 U1549 (.A1(REGISTERS[864]),
	.A2(n4008),
	.ZN(n973));
   OAI21_X1 U1550 (.A(n975),
	.B1(FE_OFN86_n4008),
	.B2(n42),
	.ZN(n1973));
   NAND2_X1 U1551 (.A1(REGISTERS[866]),
	.A2(FE_OFN86_n4008),
	.ZN(n975));
   OAI21_X1 U1552 (.A(n978),
	.B1(FE_OFN86_n4008),
	.B2(n48),
	.ZN(n1976));
   NAND2_X1 U1553 (.A1(REGISTERS[869]),
	.A2(FE_OFN86_n4008),
	.ZN(n978));
   OAI21_X1 U1554 (.A(n979),
	.B1(n4008),
	.B2(n50),
	.ZN(n1977));
   NAND2_X1 U1555 (.A1(REGISTERS[870]),
	.A2(n4008),
	.ZN(n979));
   OAI21_X1 U1556 (.A(n980),
	.B1(FE_OFN86_n4008),
	.B2(n52),
	.ZN(n1978));
   NAND2_X1 U1557 (.A1(REGISTERS[871]),
	.A2(FE_OFN86_n4008),
	.ZN(n980));
   OAI21_X1 U1558 (.A(n981),
	.B1(n4008),
	.B2(n54),
	.ZN(n1979));
   NAND2_X1 U1559 (.A1(REGISTERS[872]),
	.A2(n4008),
	.ZN(n981));
   OAI21_X1 U1560 (.A(n982),
	.B1(FE_OFN86_n4008),
	.B2(n56),
	.ZN(n1980));
   NAND2_X1 U1561 (.A1(REGISTERS[873]),
	.A2(FE_OFN86_n4008),
	.ZN(n982));
   OAI21_X1 U1562 (.A(n983),
	.B1(n4008),
	.B2(n58),
	.ZN(n1981));
   NAND2_X1 U1563 (.A1(REGISTERS[874]),
	.A2(n4008),
	.ZN(n983));
   OAI21_X1 U1564 (.A(n984),
	.B1(FE_OFN86_n4008),
	.B2(n60),
	.ZN(n1982));
   NAND2_X1 U1565 (.A1(REGISTERS[875]),
	.A2(FE_OFN86_n4008),
	.ZN(n984));
   OAI21_X1 U1566 (.A(n985),
	.B1(n4008),
	.B2(n62),
	.ZN(n1983));
   NAND2_X1 U1567 (.A1(REGISTERS[876]),
	.A2(n4008),
	.ZN(n985));
   OAI21_X1 U1568 (.A(n986),
	.B1(n4008),
	.B2(n64),
	.ZN(n1984));
   NAND2_X1 U1569 (.A1(REGISTERS[877]),
	.A2(n4008),
	.ZN(n986));
   OAI21_X1 U1570 (.A(n987),
	.B1(FE_OFN86_n4008),
	.B2(n66),
	.ZN(n1985));
   NAND2_X1 U1571 (.A1(REGISTERS[878]),
	.A2(FE_OFN86_n4008),
	.ZN(n987));
   OAI21_X1 U1572 (.A(n988),
	.B1(FE_OFN86_n4008),
	.B2(n68),
	.ZN(n1986));
   NAND2_X1 U1573 (.A1(REGISTERS[879]),
	.A2(FE_OFN86_n4008),
	.ZN(n988));
   OAI21_X1 U1574 (.A(n989),
	.B1(FE_OFN86_n4008),
	.B2(n70),
	.ZN(n1987));
   NAND2_X1 U1575 (.A1(REGISTERS[880]),
	.A2(FE_OFN86_n4008),
	.ZN(n989));
   OAI21_X1 U1576 (.A(n990),
	.B1(FE_OFN86_n4008),
	.B2(n72),
	.ZN(n1988));
   NAND2_X1 U1577 (.A1(REGISTERS[881]),
	.A2(FE_OFN86_n4008),
	.ZN(n990));
   OAI21_X1 U1578 (.A(n991),
	.B1(n4008),
	.B2(n74),
	.ZN(n1989));
   NAND2_X1 U1579 (.A1(REGISTERS[882]),
	.A2(n4008),
	.ZN(n991));
   OAI21_X1 U1580 (.A(n992),
	.B1(FE_OFN86_n4008),
	.B2(n76),
	.ZN(n1990));
   NAND2_X1 U1581 (.A1(REGISTERS[883]),
	.A2(FE_OFN86_n4008),
	.ZN(n992));
   OAI21_X1 U1582 (.A(n993),
	.B1(n4008),
	.B2(n78),
	.ZN(n1991));
   NAND2_X1 U1583 (.A1(REGISTERS[884]),
	.A2(n4008),
	.ZN(n993));
   OAI21_X1 U1584 (.A(n994),
	.B1(FE_OFN86_n4008),
	.B2(n80),
	.ZN(n1992));
   NAND2_X1 U1585 (.A1(REGISTERS[885]),
	.A2(FE_OFN86_n4008),
	.ZN(n994));
   OAI21_X1 U1586 (.A(n995),
	.B1(FE_OFN86_n4008),
	.B2(n82),
	.ZN(n1993));
   NAND2_X1 U1587 (.A1(REGISTERS[886]),
	.A2(FE_OFN86_n4008),
	.ZN(n995));
   OAI21_X1 U1588 (.A(n996),
	.B1(FE_OFN86_n4008),
	.B2(n84),
	.ZN(n1994));
   NAND2_X1 U1589 (.A1(REGISTERS[887]),
	.A2(FE_OFN86_n4008),
	.ZN(n996));
   OAI21_X1 U1590 (.A(n997),
	.B1(n4008),
	.B2(n86),
	.ZN(n1995));
   NAND2_X1 U1591 (.A1(REGISTERS[888]),
	.A2(n4008),
	.ZN(n997));
   OAI21_X1 U1592 (.A(n998),
	.B1(FE_OFN86_n4008),
	.B2(n88),
	.ZN(n1996));
   NAND2_X1 U1593 (.A1(REGISTERS[889]),
	.A2(FE_OFN86_n4008),
	.ZN(n998));
   OAI21_X1 U1594 (.A(n999),
	.B1(n4008),
	.B2(n90),
	.ZN(n1997));
   NAND2_X1 U1595 (.A1(REGISTERS[890]),
	.A2(n4008),
	.ZN(n999));
   OAI21_X1 U1596 (.A(n1000),
	.B1(FE_OFN86_n4008),
	.B2(n92),
	.ZN(n1998));
   NAND2_X1 U1597 (.A1(REGISTERS[891]),
	.A2(FE_OFN86_n4008),
	.ZN(n1000));
   OAI21_X1 U1598 (.A(n1001),
	.B1(FE_OFN86_n4008),
	.B2(n94),
	.ZN(n1999));
   NAND2_X1 U1599 (.A1(REGISTERS[892]),
	.A2(FE_OFN86_n4008),
	.ZN(n1001));
   OAI21_X1 U1600 (.A(n1006),
	.B1(n4007),
	.B2(n38),
	.ZN(n2003));
   NAND2_X1 U1601 (.A1(REGISTERS[896]),
	.A2(n4007),
	.ZN(n1006));
   OAI21_X1 U1602 (.A(n1008),
	.B1(FE_OFN82_n4007),
	.B2(n42),
	.ZN(n2005));
   NAND2_X1 U1603 (.A1(REGISTERS[898]),
	.A2(FE_OFN82_n4007),
	.ZN(n1008));
   OAI21_X1 U1604 (.A(n1011),
	.B1(FE_OFN82_n4007),
	.B2(n48),
	.ZN(n2008));
   NAND2_X1 U1605 (.A1(REGISTERS[901]),
	.A2(FE_OFN82_n4007),
	.ZN(n1011));
   OAI21_X1 U1606 (.A(n1012),
	.B1(n4007),
	.B2(n50),
	.ZN(n2009));
   NAND2_X1 U1607 (.A1(REGISTERS[902]),
	.A2(n4007),
	.ZN(n1012));
   OAI21_X1 U1608 (.A(n1013),
	.B1(FE_OFN82_n4007),
	.B2(n52),
	.ZN(n2010));
   NAND2_X1 U1609 (.A1(REGISTERS[903]),
	.A2(FE_OFN82_n4007),
	.ZN(n1013));
   OAI21_X1 U1610 (.A(n1014),
	.B1(n4007),
	.B2(n54),
	.ZN(n2011));
   NAND2_X1 U1611 (.A1(REGISTERS[904]),
	.A2(n4007),
	.ZN(n1014));
   OAI21_X1 U1612 (.A(n1015),
	.B1(FE_OFN82_n4007),
	.B2(n56),
	.ZN(n2012));
   NAND2_X1 U1613 (.A1(REGISTERS[905]),
	.A2(FE_OFN82_n4007),
	.ZN(n1015));
   OAI21_X1 U1614 (.A(n1016),
	.B1(n4007),
	.B2(n58),
	.ZN(n2013));
   NAND2_X1 U1615 (.A1(REGISTERS[906]),
	.A2(n4007),
	.ZN(n1016));
   OAI21_X1 U1616 (.A(n1017),
	.B1(FE_OFN82_n4007),
	.B2(n60),
	.ZN(n2014));
   NAND2_X1 U1617 (.A1(REGISTERS[907]),
	.A2(FE_OFN82_n4007),
	.ZN(n1017));
   OAI21_X1 U1618 (.A(n1018),
	.B1(n4007),
	.B2(n62),
	.ZN(n2015));
   NAND2_X1 U1619 (.A1(REGISTERS[908]),
	.A2(n4007),
	.ZN(n1018));
   OAI21_X1 U1620 (.A(n1019),
	.B1(n4007),
	.B2(n64),
	.ZN(n2016));
   NAND2_X1 U1621 (.A1(REGISTERS[909]),
	.A2(n4007),
	.ZN(n1019));
   OAI21_X1 U1622 (.A(n1020),
	.B1(FE_OFN82_n4007),
	.B2(n66),
	.ZN(n2017));
   NAND2_X1 U1623 (.A1(REGISTERS[910]),
	.A2(FE_OFN82_n4007),
	.ZN(n1020));
   OAI21_X1 U1624 (.A(n1021),
	.B1(FE_OFN82_n4007),
	.B2(n68),
	.ZN(n2018));
   NAND2_X1 U1625 (.A1(REGISTERS[911]),
	.A2(FE_OFN82_n4007),
	.ZN(n1021));
   OAI21_X1 U1626 (.A(n1022),
	.B1(FE_OFN82_n4007),
	.B2(n70),
	.ZN(n2019));
   NAND2_X1 U1627 (.A1(REGISTERS[912]),
	.A2(FE_OFN82_n4007),
	.ZN(n1022));
   OAI21_X1 U1628 (.A(n1023),
	.B1(FE_OFN82_n4007),
	.B2(n72),
	.ZN(n2020));
   NAND2_X1 U1629 (.A1(REGISTERS[913]),
	.A2(FE_OFN82_n4007),
	.ZN(n1023));
   OAI21_X1 U1630 (.A(n1024),
	.B1(n4007),
	.B2(n74),
	.ZN(n2021));
   NAND2_X1 U1631 (.A1(REGISTERS[914]),
	.A2(n4007),
	.ZN(n1024));
   OAI21_X1 U1632 (.A(n1025),
	.B1(FE_OFN82_n4007),
	.B2(n76),
	.ZN(n2022));
   NAND2_X1 U1633 (.A1(REGISTERS[915]),
	.A2(FE_OFN82_n4007),
	.ZN(n1025));
   OAI21_X1 U1634 (.A(n1026),
	.B1(n4007),
	.B2(n78),
	.ZN(n2023));
   NAND2_X1 U1635 (.A1(REGISTERS[916]),
	.A2(n4007),
	.ZN(n1026));
   OAI21_X1 U1636 (.A(n1027),
	.B1(FE_OFN82_n4007),
	.B2(n80),
	.ZN(n2024));
   NAND2_X1 U1637 (.A1(REGISTERS[917]),
	.A2(FE_OFN82_n4007),
	.ZN(n1027));
   OAI21_X1 U1638 (.A(n1028),
	.B1(FE_OFN82_n4007),
	.B2(n82),
	.ZN(n2025));
   NAND2_X1 U1639 (.A1(REGISTERS[918]),
	.A2(FE_OFN82_n4007),
	.ZN(n1028));
   OAI21_X1 U1640 (.A(n1029),
	.B1(FE_OFN82_n4007),
	.B2(n84),
	.ZN(n2026));
   NAND2_X1 U1641 (.A1(REGISTERS[919]),
	.A2(FE_OFN82_n4007),
	.ZN(n1029));
   OAI21_X1 U1642 (.A(n1030),
	.B1(n4007),
	.B2(n86),
	.ZN(n2027));
   NAND2_X1 U1643 (.A1(REGISTERS[920]),
	.A2(n4007),
	.ZN(n1030));
   OAI21_X1 U1644 (.A(n1031),
	.B1(FE_OFN82_n4007),
	.B2(n88),
	.ZN(n2028));
   NAND2_X1 U1645 (.A1(REGISTERS[921]),
	.A2(FE_OFN82_n4007),
	.ZN(n1031));
   OAI21_X1 U1646 (.A(n1032),
	.B1(n4007),
	.B2(n90),
	.ZN(n2029));
   NAND2_X1 U1647 (.A1(REGISTERS[922]),
	.A2(n4007),
	.ZN(n1032));
   OAI21_X1 U1648 (.A(n1033),
	.B1(FE_OFN82_n4007),
	.B2(n92),
	.ZN(n2030));
   NAND2_X1 U1649 (.A1(REGISTERS[923]),
	.A2(FE_OFN82_n4007),
	.ZN(n1033));
   OAI21_X1 U1650 (.A(n1034),
	.B1(FE_OFN82_n4007),
	.B2(n94),
	.ZN(n2031));
   NAND2_X1 U1651 (.A1(REGISTERS[924]),
	.A2(FE_OFN82_n4007),
	.ZN(n1034));
   OAI21_X1 U1652 (.A(n1039),
	.B1(FE_OFN71_n4006),
	.B2(n38),
	.ZN(n2035));
   NAND2_X1 U1653 (.A1(REGISTERS[928]),
	.A2(FE_OFN71_n4006),
	.ZN(n1039));
   OAI21_X1 U1654 (.A(n1041),
	.B1(FE_OFN71_n4006),
	.B2(n42),
	.ZN(n2037));
   NAND2_X1 U1655 (.A1(REGISTERS[930]),
	.A2(FE_OFN71_n4006),
	.ZN(n1041));
   OAI21_X1 U1656 (.A(n1044),
	.B1(FE_OFN71_n4006),
	.B2(n48),
	.ZN(n2040));
   NAND2_X1 U1657 (.A1(REGISTERS[933]),
	.A2(FE_OFN71_n4006),
	.ZN(n1044));
   OAI21_X1 U1658 (.A(n1045),
	.B1(FE_OFN71_n4006),
	.B2(n50),
	.ZN(n2041));
   NAND2_X1 U1659 (.A1(REGISTERS[934]),
	.A2(FE_OFN71_n4006),
	.ZN(n1045));
   OAI21_X1 U1660 (.A(n1046),
	.B1(FE_OFN71_n4006),
	.B2(n52),
	.ZN(n2042));
   NAND2_X1 U1661 (.A1(REGISTERS[935]),
	.A2(FE_OFN71_n4006),
	.ZN(n1046));
   OAI21_X1 U1662 (.A(n1047),
	.B1(FE_OFN71_n4006),
	.B2(n54),
	.ZN(n2043));
   NAND2_X1 U1663 (.A1(REGISTERS[936]),
	.A2(FE_OFN71_n4006),
	.ZN(n1047));
   OAI21_X1 U1664 (.A(n1048),
	.B1(n4006),
	.B2(n56),
	.ZN(n2044));
   NAND2_X1 U1665 (.A1(REGISTERS[937]),
	.A2(n4006),
	.ZN(n1048));
   OAI21_X1 U1666 (.A(n1049),
	.B1(FE_OFN71_n4006),
	.B2(n58),
	.ZN(n2045));
   NAND2_X1 U1667 (.A1(REGISTERS[938]),
	.A2(FE_OFN71_n4006),
	.ZN(n1049));
   OAI21_X1 U1668 (.A(n1050),
	.B1(n4006),
	.B2(n60),
	.ZN(n2046));
   NAND2_X1 U1669 (.A1(REGISTERS[939]),
	.A2(n4006),
	.ZN(n1050));
   OAI21_X1 U1670 (.A(n1051),
	.B1(FE_OFN71_n4006),
	.B2(n62),
	.ZN(n2047));
   NAND2_X1 U1671 (.A1(REGISTERS[940]),
	.A2(FE_OFN71_n4006),
	.ZN(n1051));
   OAI21_X1 U1672 (.A(n1052),
	.B1(FE_OFN71_n4006),
	.B2(n64),
	.ZN(n2048));
   NAND2_X1 U1673 (.A1(REGISTERS[941]),
	.A2(FE_OFN71_n4006),
	.ZN(n1052));
   OAI21_X1 U1674 (.A(n1053),
	.B1(FE_OFN71_n4006),
	.B2(n66),
	.ZN(n2049));
   NAND2_X1 U1675 (.A1(REGISTERS[942]),
	.A2(FE_OFN71_n4006),
	.ZN(n1053));
   OAI21_X1 U1676 (.A(n1054),
	.B1(FE_OFN71_n4006),
	.B2(n68),
	.ZN(n2050));
   NAND2_X1 U1677 (.A1(REGISTERS[943]),
	.A2(FE_OFN71_n4006),
	.ZN(n1054));
   OAI21_X1 U1678 (.A(n1055),
	.B1(n4006),
	.B2(n70),
	.ZN(n2051));
   NAND2_X1 U1679 (.A1(REGISTERS[944]),
	.A2(n4006),
	.ZN(n1055));
   OAI21_X1 U1680 (.A(n1056),
	.B1(FE_OFN71_n4006),
	.B2(n72),
	.ZN(n2052));
   NAND2_X1 U1681 (.A1(REGISTERS[945]),
	.A2(FE_OFN71_n4006),
	.ZN(n1056));
   OAI21_X1 U1682 (.A(n1057),
	.B1(FE_OFN71_n4006),
	.B2(n74),
	.ZN(n2053));
   NAND2_X1 U1683 (.A1(REGISTERS[946]),
	.A2(FE_OFN71_n4006),
	.ZN(n1057));
   OAI21_X1 U1684 (.A(n1058),
	.B1(FE_OFN71_n4006),
	.B2(n76),
	.ZN(n2054));
   NAND2_X1 U1685 (.A1(REGISTERS[947]),
	.A2(FE_OFN71_n4006),
	.ZN(n1058));
   OAI21_X1 U1686 (.A(n1059),
	.B1(FE_OFN71_n4006),
	.B2(n78),
	.ZN(n2055));
   NAND2_X1 U1687 (.A1(REGISTERS[948]),
	.A2(FE_OFN71_n4006),
	.ZN(n1059));
   OAI21_X1 U1688 (.A(n1060),
	.B1(FE_OFN71_n4006),
	.B2(n80),
	.ZN(n2056));
   NAND2_X1 U1689 (.A1(REGISTERS[949]),
	.A2(FE_OFN71_n4006),
	.ZN(n1060));
   OAI21_X1 U1690 (.A(n1061),
	.B1(FE_OFN71_n4006),
	.B2(n82),
	.ZN(n2057));
   NAND2_X1 U1691 (.A1(REGISTERS[950]),
	.A2(FE_OFN71_n4006),
	.ZN(n1061));
   OAI21_X1 U1692 (.A(n1062),
	.B1(FE_OFN71_n4006),
	.B2(n84),
	.ZN(n2058));
   NAND2_X1 U1693 (.A1(REGISTERS[951]),
	.A2(FE_OFN71_n4006),
	.ZN(n1062));
   OAI21_X1 U1694 (.A(n1063),
	.B1(FE_OFN71_n4006),
	.B2(n86),
	.ZN(n2059));
   NAND2_X1 U1695 (.A1(REGISTERS[952]),
	.A2(FE_OFN71_n4006),
	.ZN(n1063));
   OAI21_X1 U1696 (.A(n1064),
	.B1(FE_OFN71_n4006),
	.B2(n88),
	.ZN(n2060));
   NAND2_X1 U1697 (.A1(REGISTERS[953]),
	.A2(FE_OFN71_n4006),
	.ZN(n1064));
   OAI21_X1 U1698 (.A(n1065),
	.B1(FE_OFN71_n4006),
	.B2(n90),
	.ZN(n2061));
   NAND2_X1 U1699 (.A1(REGISTERS[954]),
	.A2(FE_OFN71_n4006),
	.ZN(n1065));
   OAI21_X1 U1700 (.A(n1066),
	.B1(FE_OFN71_n4006),
	.B2(n92),
	.ZN(n2062));
   NAND2_X1 U1701 (.A1(REGISTERS[955]),
	.A2(FE_OFN71_n4006),
	.ZN(n1066));
   OAI21_X1 U1702 (.A(n1067),
	.B1(FE_OFN71_n4006),
	.B2(n94),
	.ZN(n2063));
   NAND2_X1 U1703 (.A1(REGISTERS[956]),
	.A2(FE_OFN71_n4006),
	.ZN(n1067));
   OAI21_X1 U1704 (.A(n1079),
	.B1(FE_OFN84_n4005),
	.B2(n52),
	.ZN(n2074));
   NAND2_X1 U1705 (.A1(REGISTERS[967]),
	.A2(FE_OFN84_n4005),
	.ZN(n1079));
   OAI21_X1 U1706 (.A(n1080),
	.B1(n4005),
	.B2(n54),
	.ZN(n2075));
   NAND2_X1 U1707 (.A1(REGISTERS[968]),
	.A2(n4005),
	.ZN(n1080));
   OAI21_X1 U1708 (.A(n1081),
	.B1(FE_OFN84_n4005),
	.B2(n56),
	.ZN(n2076));
   NAND2_X1 U1709 (.A1(REGISTERS[969]),
	.A2(FE_OFN84_n4005),
	.ZN(n1081));
   OAI21_X1 U1710 (.A(n1082),
	.B1(n4005),
	.B2(n58),
	.ZN(n2077));
   NAND2_X1 U1711 (.A1(REGISTERS[970]),
	.A2(n4005),
	.ZN(n1082));
   OAI21_X1 U1712 (.A(n1083),
	.B1(FE_OFN84_n4005),
	.B2(n60),
	.ZN(n2078));
   NAND2_X1 U1713 (.A1(REGISTERS[971]),
	.A2(FE_OFN84_n4005),
	.ZN(n1083));
   OAI21_X1 U1714 (.A(n1084),
	.B1(n4005),
	.B2(n62),
	.ZN(n2079));
   NAND2_X1 U1715 (.A1(REGISTERS[972]),
	.A2(n4005),
	.ZN(n1084));
   OAI21_X1 U1716 (.A(n1086),
	.B1(FE_OFN84_n4005),
	.B2(n66),
	.ZN(n2081));
   NAND2_X1 U1717 (.A1(REGISTERS[974]),
	.A2(FE_OFN84_n4005),
	.ZN(n1086));
   OAI21_X1 U1718 (.A(n1087),
	.B1(FE_OFN84_n4005),
	.B2(n68),
	.ZN(n2082));
   NAND2_X1 U1719 (.A1(REGISTERS[975]),
	.A2(FE_OFN84_n4005),
	.ZN(n1087));
   OAI21_X1 U1720 (.A(n208),
	.B1(n4024),
	.B2(n40),
	.ZN(n1236));
   NAND2_X1 U1721 (.A1(REGISTERS[129]),
	.A2(n4024),
	.ZN(n208));
   OAI21_X1 U1722 (.A(n210),
	.B1(FE_OFN83_n4024),
	.B2(n44),
	.ZN(n1238));
   NAND2_X1 U1723 (.A1(REGISTERS[131]),
	.A2(FE_OFN83_n4024),
	.ZN(n210));
   OAI21_X1 U1724 (.A(n211),
	.B1(n4024),
	.B2(n46),
	.ZN(n1239));
   NAND2_X1 U1725 (.A1(REGISTERS[132]),
	.A2(n4024),
	.ZN(n211));
   OAI21_X1 U1726 (.A(n238),
	.B1(n4024),
	.B2(n100),
	.ZN(n1266));
   NAND2_X1 U1727 (.A1(REGISTERS[159]),
	.A2(n4024),
	.ZN(n238));
   OAI21_X1 U1728 (.A(n344),
	.B1(n4036),
	.B2(n40),
	.ZN(n1364));
   NAND2_X1 U1729 (.A1(REGISTERS[257]),
	.A2(n4036),
	.ZN(n344));
   OAI21_X1 U1730 (.A(n346),
	.B1(FE_OFN60_n4036),
	.B2(n44),
	.ZN(n1366));
   NAND2_X1 U1731 (.A1(REGISTERS[259]),
	.A2(FE_OFN60_n4036),
	.ZN(n346));
   OAI21_X1 U1732 (.A(n347),
	.B1(n4036),
	.B2(n46),
	.ZN(n1367));
   NAND2_X1 U1733 (.A1(REGISTERS[260]),
	.A2(n4036),
	.ZN(n347));
   OAI21_X1 U1734 (.A(n374),
	.B1(n4036),
	.B2(n100),
	.ZN(n1394));
   NAND2_X1 U1735 (.A1(REGISTERS[287]),
	.A2(n4036),
	.ZN(n374));
   OAI21_X1 U1736 (.A(n378),
	.B1(n4035),
	.B2(n40),
	.ZN(n1396));
   NAND2_X1 U1737 (.A1(REGISTERS[289]),
	.A2(n4035),
	.ZN(n378));
   OAI21_X1 U1738 (.A(n380),
	.B1(FE_OFN80_n4035),
	.B2(n44),
	.ZN(n1398));
   NAND2_X1 U1739 (.A1(REGISTERS[291]),
	.A2(FE_OFN80_n4035),
	.ZN(n380));
   OAI21_X1 U1740 (.A(n381),
	.B1(n4035),
	.B2(n46),
	.ZN(n1399));
   NAND2_X1 U1741 (.A1(REGISTERS[292]),
	.A2(n4035),
	.ZN(n381));
   OAI21_X1 U1742 (.A(n408),
	.B1(n4035),
	.B2(n100),
	.ZN(n1426));
   NAND2_X1 U1743 (.A1(REGISTERS[319]),
	.A2(n4035),
	.ZN(n408));
   OAI21_X1 U1744 (.A(n411),
	.B1(FE_OFN59_n4034),
	.B2(n40),
	.ZN(n1428));
   NAND2_X1 U1745 (.A1(REGISTERS[321]),
	.A2(FE_OFN59_n4034),
	.ZN(n411));
   OAI21_X1 U1746 (.A(n413),
	.B1(FE_OFN59_n4034),
	.B2(n44),
	.ZN(n1430));
   NAND2_X1 U1747 (.A1(REGISTERS[323]),
	.A2(FE_OFN59_n4034),
	.ZN(n413));
   OAI21_X1 U1748 (.A(n414),
	.B1(n4034),
	.B2(n46),
	.ZN(n1431));
   NAND2_X1 U1749 (.A1(REGISTERS[324]),
	.A2(n4034),
	.ZN(n414));
   OAI21_X1 U1750 (.A(n441),
	.B1(FE_OFN59_n4034),
	.B2(n100),
	.ZN(n1458));
   NAND2_X1 U1751 (.A1(REGISTERS[351]),
	.A2(FE_OFN59_n4034),
	.ZN(n441));
   OAI21_X1 U1752 (.A(n444),
	.B1(FE_OFN70_n4033),
	.B2(n40),
	.ZN(n1460));
   NAND2_X1 U1753 (.A1(REGISTERS[353]),
	.A2(FE_OFN70_n4033),
	.ZN(n444));
   OAI21_X1 U1754 (.A(n446),
	.B1(FE_OFN70_n4033),
	.B2(n44),
	.ZN(n1462));
   NAND2_X1 U1755 (.A1(REGISTERS[355]),
	.A2(FE_OFN70_n4033),
	.ZN(n446));
   OAI21_X1 U1756 (.A(n447),
	.B1(n4033),
	.B2(n46),
	.ZN(n1463));
   NAND2_X1 U1757 (.A1(REGISTERS[356]),
	.A2(n4033),
	.ZN(n447));
   OAI21_X1 U1758 (.A(n474),
	.B1(FE_OFN70_n4033),
	.B2(n100),
	.ZN(n1490));
   NAND2_X1 U1759 (.A1(REGISTERS[383]),
	.A2(FE_OFN70_n4033),
	.ZN(n474));
   OAI21_X1 U1760 (.A(n477),
	.B1(n4032),
	.B2(n40),
	.ZN(n1492));
   NAND2_X1 U1761 (.A1(REGISTERS[385]),
	.A2(n4032),
	.ZN(n477));
   OAI21_X1 U1762 (.A(n479),
	.B1(FE_OFN87_n4032),
	.B2(n44),
	.ZN(n1494));
   NAND2_X1 U1763 (.A1(REGISTERS[387]),
	.A2(FE_OFN87_n4032),
	.ZN(n479));
   OAI21_X1 U1764 (.A(n480),
	.B1(n4032),
	.B2(n46),
	.ZN(n1495));
   NAND2_X1 U1765 (.A1(REGISTERS[388]),
	.A2(n4032),
	.ZN(n480));
   OAI21_X1 U1766 (.A(n507),
	.B1(n4032),
	.B2(n100),
	.ZN(n1522));
   NAND2_X1 U1767 (.A1(REGISTERS[415]),
	.A2(n4032),
	.ZN(n507));
   OAI21_X1 U1768 (.A(n510),
	.B1(FE_OFN63_n4031),
	.B2(n40),
	.ZN(n1524));
   NAND2_X1 U1769 (.A1(REGISTERS[417]),
	.A2(FE_OFN63_n4031),
	.ZN(n510));
   OAI21_X1 U1770 (.A(n512),
	.B1(FE_OFN63_n4031),
	.B2(n44),
	.ZN(n1526));
   NAND2_X1 U1771 (.A1(REGISTERS[419]),
	.A2(FE_OFN63_n4031),
	.ZN(n512));
   OAI21_X1 U1772 (.A(n513),
	.B1(n4031),
	.B2(n46),
	.ZN(n1527));
   NAND2_X1 U1773 (.A1(REGISTERS[420]),
	.A2(n4031),
	.ZN(n513));
   OAI21_X1 U1774 (.A(n540),
	.B1(FE_OFN63_n4031),
	.B2(n100),
	.ZN(n1554));
   NAND2_X1 U1775 (.A1(REGISTERS[447]),
	.A2(FE_OFN63_n4031),
	.ZN(n540));
   OAI21_X1 U1776 (.A(n543),
	.B1(n4030),
	.B2(n40),
	.ZN(n1556));
   NAND2_X1 U1777 (.A1(REGISTERS[449]),
	.A2(n4030),
	.ZN(n543));
   OAI21_X1 U1778 (.A(n545),
	.B1(FE_OFN81_n4030),
	.B2(n44),
	.ZN(n1558));
   NAND2_X1 U1779 (.A1(REGISTERS[451]),
	.A2(FE_OFN81_n4030),
	.ZN(n545));
   OAI21_X1 U1780 (.A(n546),
	.B1(n4030),
	.B2(n46),
	.ZN(n1559));
   NAND2_X1 U1781 (.A1(REGISTERS[452]),
	.A2(n4030),
	.ZN(n546));
   OAI21_X1 U1782 (.A(n573),
	.B1(n4030),
	.B2(n100),
	.ZN(n1586));
   NAND2_X1 U1783 (.A1(REGISTERS[479]),
	.A2(n4030),
	.ZN(n573));
   OAI21_X1 U1784 (.A(n576),
	.B1(n4029),
	.B2(n40),
	.ZN(n1588));
   NAND2_X1 U1785 (.A1(REGISTERS[481]),
	.A2(n4029),
	.ZN(n576));
   OAI21_X1 U1786 (.A(n578),
	.B1(FE_OFN67_n4029),
	.B2(n44),
	.ZN(n1590));
   NAND2_X1 U1787 (.A1(REGISTERS[483]),
	.A2(FE_OFN67_n4029),
	.ZN(n578));
   OAI21_X1 U1788 (.A(n579),
	.B1(n4029),
	.B2(n46),
	.ZN(n1591));
   NAND2_X1 U1789 (.A1(REGISTERS[484]),
	.A2(n4029),
	.ZN(n579));
   OAI21_X1 U1790 (.A(n606),
	.B1(n4029),
	.B2(n100),
	.ZN(n1618));
   NAND2_X1 U1791 (.A1(REGISTERS[511]),
	.A2(n4029),
	.ZN(n606));
   OAI21_X1 U1792 (.A(n609),
	.B1(n4019),
	.B2(n40),
	.ZN(n1620));
   NAND2_X1 U1793 (.A1(REGISTERS[513]),
	.A2(n4019),
	.ZN(n609));
   OAI21_X1 U1794 (.A(n611),
	.B1(FE_OFN61_n4019),
	.B2(n44),
	.ZN(n1622));
   NAND2_X1 U1795 (.A1(REGISTERS[515]),
	.A2(FE_OFN61_n4019),
	.ZN(n611));
   OAI21_X1 U1796 (.A(n612),
	.B1(n4019),
	.B2(n46),
	.ZN(n1623));
   NAND2_X1 U1797 (.A1(REGISTERS[516]),
	.A2(n4019),
	.ZN(n612));
   OAI21_X1 U1798 (.A(n639),
	.B1(FE_OFN61_n4019),
	.B2(n100),
	.ZN(n1650));
   NAND2_X1 U1799 (.A1(REGISTERS[543]),
	.A2(FE_OFN61_n4019),
	.ZN(n639));
   OAI21_X1 U1800 (.A(n643),
	.B1(FE_OFN65_n4018),
	.B2(n40),
	.ZN(n1652));
   NAND2_X1 U1801 (.A1(REGISTERS[545]),
	.A2(FE_OFN65_n4018),
	.ZN(n643));
   OAI21_X1 U1802 (.A(n645),
	.B1(FE_OFN65_n4018),
	.B2(n44),
	.ZN(n1654));
   NAND2_X1 U1803 (.A1(REGISTERS[547]),
	.A2(FE_OFN65_n4018),
	.ZN(n645));
   OAI21_X1 U1804 (.A(n646),
	.B1(n4018),
	.B2(n46),
	.ZN(n1655));
   NAND2_X1 U1805 (.A1(REGISTERS[548]),
	.A2(n4018),
	.ZN(n646));
   OAI21_X1 U1806 (.A(n673),
	.B1(FE_OFN65_n4018),
	.B2(n100),
	.ZN(n1682));
   NAND2_X1 U1807 (.A1(REGISTERS[575]),
	.A2(FE_OFN65_n4018),
	.ZN(n673));
   OAI21_X1 U1808 (.A(n676),
	.B1(n4017),
	.B2(n40),
	.ZN(n1684));
   NAND2_X1 U1809 (.A1(REGISTERS[577]),
	.A2(n4017),
	.ZN(n676));
   OAI21_X1 U1810 (.A(n678),
	.B1(FE_OFN66_n4017),
	.B2(n44),
	.ZN(n1686));
   NAND2_X1 U1811 (.A1(REGISTERS[579]),
	.A2(FE_OFN66_n4017),
	.ZN(n678));
   OAI21_X1 U1812 (.A(n679),
	.B1(FE_OFN66_n4017),
	.B2(n46),
	.ZN(n1687));
   NAND2_X1 U1813 (.A1(REGISTERS[580]),
	.A2(FE_OFN66_n4017),
	.ZN(n679));
   OAI21_X1 U1814 (.A(n706),
	.B1(FE_OFN66_n4017),
	.B2(n100),
	.ZN(n1714));
   NAND2_X1 U1815 (.A1(REGISTERS[607]),
	.A2(FE_OFN66_n4017),
	.ZN(n706));
   OAI21_X1 U1816 (.A(n709),
	.B1(FE_OFN62_n4016),
	.B2(n40),
	.ZN(n1716));
   NAND2_X1 U1817 (.A1(REGISTERS[609]),
	.A2(FE_OFN62_n4016),
	.ZN(n709));
   OAI21_X1 U1818 (.A(n711),
	.B1(FE_OFN62_n4016),
	.B2(n44),
	.ZN(n1718));
   NAND2_X1 U1819 (.A1(REGISTERS[611]),
	.A2(FE_OFN62_n4016),
	.ZN(n711));
   OAI21_X1 U1820 (.A(n712),
	.B1(n4016),
	.B2(n46),
	.ZN(n1719));
   NAND2_X1 U1821 (.A1(REGISTERS[612]),
	.A2(n4016),
	.ZN(n712));
   OAI21_X1 U1822 (.A(n739),
	.B1(FE_OFN62_n4016),
	.B2(n100),
	.ZN(n1746));
   NAND2_X1 U1823 (.A1(REGISTERS[639]),
	.A2(FE_OFN62_n4016),
	.ZN(n739));
   OAI21_X1 U1824 (.A(n742),
	.B1(n4015),
	.B2(n40),
	.ZN(n1748));
   NAND2_X1 U1825 (.A1(REGISTERS[641]),
	.A2(n4015),
	.ZN(n742));
   OAI21_X1 U1826 (.A(n744),
	.B1(FE_OFN74_n4015),
	.B2(n44),
	.ZN(n1750));
   NAND2_X1 U1827 (.A1(REGISTERS[643]),
	.A2(FE_OFN74_n4015),
	.ZN(n744));
   OAI21_X1 U1828 (.A(n745),
	.B1(n4015),
	.B2(n46),
	.ZN(n1751));
   NAND2_X1 U1829 (.A1(REGISTERS[644]),
	.A2(n4015),
	.ZN(n745));
   OAI21_X1 U1830 (.A(n772),
	.B1(n4015),
	.B2(n100),
	.ZN(n1778));
   NAND2_X1 U1831 (.A1(REGISTERS[671]),
	.A2(n4015),
	.ZN(n772));
   OAI21_X1 U1832 (.A(n775),
	.B1(n4014),
	.B2(n40),
	.ZN(n1780));
   NAND2_X1 U1833 (.A1(REGISTERS[673]),
	.A2(n4014),
	.ZN(n775));
   OAI21_X1 U1834 (.A(n777),
	.B1(FE_OFN78_n4014),
	.B2(n44),
	.ZN(n1782));
   NAND2_X1 U1835 (.A1(REGISTERS[675]),
	.A2(FE_OFN78_n4014),
	.ZN(n777));
   OAI21_X1 U1836 (.A(n778),
	.B1(n4014),
	.B2(n46),
	.ZN(n1783));
   NAND2_X1 U1837 (.A1(REGISTERS[676]),
	.A2(n4014),
	.ZN(n778));
   OAI21_X1 U1838 (.A(n805),
	.B1(FE_OFN78_n4014),
	.B2(n100),
	.ZN(n1810));
   NAND2_X1 U1839 (.A1(REGISTERS[703]),
	.A2(FE_OFN78_n4014),
	.ZN(n805));
   OAI21_X1 U1840 (.A(n808),
	.B1(n4013),
	.B2(n40),
	.ZN(n1812));
   NAND2_X1 U1841 (.A1(REGISTERS[705]),
	.A2(n4013),
	.ZN(n808));
   OAI21_X1 U1842 (.A(n810),
	.B1(FE_OFN76_n4013),
	.B2(n44),
	.ZN(n1814));
   NAND2_X1 U1843 (.A1(REGISTERS[707]),
	.A2(FE_OFN76_n4013),
	.ZN(n810));
   OAI21_X1 U1844 (.A(n811),
	.B1(n4013),
	.B2(n46),
	.ZN(n1815));
   NAND2_X1 U1845 (.A1(REGISTERS[708]),
	.A2(n4013),
	.ZN(n811));
   OAI21_X1 U1846 (.A(n838),
	.B1(n4013),
	.B2(n100),
	.ZN(n1842));
   NAND2_X1 U1847 (.A1(REGISTERS[735]),
	.A2(n4013),
	.ZN(n838));
   OAI21_X1 U1848 (.A(n841),
	.B1(n4012),
	.B2(n40),
	.ZN(n1844));
   NAND2_X1 U1849 (.A1(REGISTERS[737]),
	.A2(n4012),
	.ZN(n841));
   OAI21_X1 U1850 (.A(n843),
	.B1(FE_OFN64_n4012),
	.B2(n44),
	.ZN(n1846));
   NAND2_X1 U1851 (.A1(REGISTERS[739]),
	.A2(FE_OFN64_n4012),
	.ZN(n843));
   OAI21_X1 U1852 (.A(n844),
	.B1(n4012),
	.B2(n46),
	.ZN(n1847));
   NAND2_X1 U1853 (.A1(REGISTERS[740]),
	.A2(n4012),
	.ZN(n844));
   OAI21_X1 U1854 (.A(n871),
	.B1(FE_OFN64_n4012),
	.B2(n100),
	.ZN(n1874));
   NAND2_X1 U1855 (.A1(REGISTERS[767]),
	.A2(FE_OFN64_n4012),
	.ZN(n871));
   OAI21_X1 U1856 (.A(n874),
	.B1(n4011),
	.B2(n40),
	.ZN(n1876));
   NAND2_X1 U1857 (.A1(REGISTERS[769]),
	.A2(n4011),
	.ZN(n874));
   OAI21_X1 U1858 (.A(n876),
	.B1(FE_OFN68_n4011),
	.B2(n44),
	.ZN(n1878));
   NAND2_X1 U1859 (.A1(REGISTERS[771]),
	.A2(FE_OFN68_n4011),
	.ZN(n876));
   OAI21_X1 U1860 (.A(n877),
	.B1(n4011),
	.B2(n46),
	.ZN(n1879));
   NAND2_X1 U1861 (.A1(REGISTERS[772]),
	.A2(n4011),
	.ZN(n877));
   OAI21_X1 U1862 (.A(n904),
	.B1(n4011),
	.B2(n100),
	.ZN(n1906));
   NAND2_X1 U1863 (.A1(REGISTERS[799]),
	.A2(n4011),
	.ZN(n904));
   OAI21_X1 U1864 (.A(n908),
	.B1(n4010),
	.B2(n40),
	.ZN(n1908));
   NAND2_X1 U1865 (.A1(REGISTERS[801]),
	.A2(n4010),
	.ZN(n908));
   OAI21_X1 U1866 (.A(n910),
	.B1(FE_OFN88_n4010),
	.B2(n44),
	.ZN(n1910));
   NAND2_X1 U1867 (.A1(REGISTERS[803]),
	.A2(FE_OFN88_n4010),
	.ZN(n910));
   OAI21_X1 U1868 (.A(n911),
	.B1(FE_OFN88_n4010),
	.B2(n46),
	.ZN(n1911));
   NAND2_X1 U1869 (.A1(REGISTERS[804]),
	.A2(FE_OFN88_n4010),
	.ZN(n911));
   OAI21_X1 U1870 (.A(n938),
	.B1(n4010),
	.B2(n100),
	.ZN(n1938));
   NAND2_X1 U1871 (.A1(REGISTERS[831]),
	.A2(n4010),
	.ZN(n938));
   OAI21_X1 U1872 (.A(n941),
	.B1(n4009),
	.B2(n40),
	.ZN(n1940));
   NAND2_X1 U1873 (.A1(REGISTERS[833]),
	.A2(n4009),
	.ZN(n941));
   OAI21_X1 U1874 (.A(n943),
	.B1(FE_OFN73_n4009),
	.B2(n44),
	.ZN(n1942));
   NAND2_X1 U1875 (.A1(REGISTERS[835]),
	.A2(FE_OFN73_n4009),
	.ZN(n943));
   OAI21_X1 U1876 (.A(n944),
	.B1(FE_OFN73_n4009),
	.B2(n46),
	.ZN(n1943));
   NAND2_X1 U1877 (.A1(REGISTERS[836]),
	.A2(n4009),
	.ZN(n944));
   OAI21_X1 U1878 (.A(n971),
	.B1(n4009),
	.B2(n100),
	.ZN(n1970));
   NAND2_X1 U1879 (.A1(REGISTERS[863]),
	.A2(n4009),
	.ZN(n971));
   OAI21_X1 U1880 (.A(n974),
	.B1(n4008),
	.B2(n40),
	.ZN(n1972));
   NAND2_X1 U1881 (.A1(REGISTERS[865]),
	.A2(n4008),
	.ZN(n974));
   OAI21_X1 U1882 (.A(n976),
	.B1(FE_OFN86_n4008),
	.B2(n44),
	.ZN(n1974));
   NAND2_X1 U1883 (.A1(REGISTERS[867]),
	.A2(FE_OFN86_n4008),
	.ZN(n976));
   OAI21_X1 U1884 (.A(n977),
	.B1(FE_OFN86_n4008),
	.B2(n46),
	.ZN(n1975));
   NAND2_X1 U1885 (.A1(REGISTERS[868]),
	.A2(FE_OFN86_n4008),
	.ZN(n977));
   OAI21_X1 U1886 (.A(n1004),
	.B1(n4008),
	.B2(n100),
	.ZN(n2002));
   NAND2_X1 U1887 (.A1(REGISTERS[895]),
	.A2(n4008),
	.ZN(n1004));
   OAI21_X1 U1888 (.A(n1007),
	.B1(n4007),
	.B2(n40),
	.ZN(n2004));
   NAND2_X1 U1889 (.A1(REGISTERS[897]),
	.A2(n4007),
	.ZN(n1007));
   OAI21_X1 U1890 (.A(n1009),
	.B1(FE_OFN82_n4007),
	.B2(n44),
	.ZN(n2006));
   NAND2_X1 U1891 (.A1(REGISTERS[899]),
	.A2(FE_OFN82_n4007),
	.ZN(n1009));
   OAI21_X1 U1892 (.A(n1010),
	.B1(FE_OFN82_n4007),
	.B2(n46),
	.ZN(n2007));
   NAND2_X1 U1893 (.A1(REGISTERS[900]),
	.A2(FE_OFN82_n4007),
	.ZN(n1010));
   OAI21_X1 U1894 (.A(n1037),
	.B1(n4007),
	.B2(n100),
	.ZN(n2034));
   NAND2_X1 U1895 (.A1(REGISTERS[927]),
	.A2(n4007),
	.ZN(n1037));
   OAI21_X1 U1896 (.A(n1040),
	.B1(FE_OFN71_n4006),
	.B2(n40),
	.ZN(n2036));
   NAND2_X1 U1897 (.A1(REGISTERS[929]),
	.A2(FE_OFN71_n4006),
	.ZN(n1040));
   OAI21_X1 U1898 (.A(n1042),
	.B1(FE_OFN71_n4006),
	.B2(n44),
	.ZN(n2038));
   NAND2_X1 U1899 (.A1(REGISTERS[931]),
	.A2(FE_OFN71_n4006),
	.ZN(n1042));
   OAI21_X1 U1900 (.A(n1043),
	.B1(n4006),
	.B2(n46),
	.ZN(n2039));
   NAND2_X1 U1901 (.A1(REGISTERS[932]),
	.A2(n4006),
	.ZN(n1043));
   OAI21_X1 U1902 (.A(n1070),
	.B1(FE_OFN71_n4006),
	.B2(n100),
	.ZN(n2066));
   NAND2_X1 U1903 (.A1(REGISTERS[959]),
	.A2(FE_OFN71_n4006),
	.ZN(n1070));
   INV_X4 U1904 (.A(RESET),
	.ZN(n4041));
   INV_X1 U1905 (.A(ADD_WR[1]),
	.ZN(n4039));
   INV_X1 U1906 (.A(ADD_WR[3]),
	.ZN(n4037));
   INV_X1 U1907 (.A(ADD_WR[4]),
	.ZN(n4020));
   OAI21_X1 U1908 (.A(n236),
	.B1(FE_OFN83_n4024),
	.B2(n96),
	.ZN(n1264));
   NAND2_X1 U1909 (.A1(REGISTERS[157]),
	.A2(FE_OFN83_n4024),
	.ZN(n236));
   OAI21_X1 U1910 (.A(n237),
	.B1(FE_OFN83_n4024),
	.B2(n98),
	.ZN(n1265));
   NAND2_X1 U1911 (.A1(REGISTERS[158]),
	.A2(FE_OFN83_n4024),
	.ZN(n237));
   OAI21_X1 U1912 (.A(n350),
	.B1(FE_OFN60_n4036),
	.B2(n52),
	.ZN(n1370));
   NAND2_X1 U1913 (.A1(REGISTERS[263]),
	.A2(FE_OFN60_n4036),
	.ZN(n350));
   OAI21_X1 U1914 (.A(n351),
	.B1(n4036),
	.B2(n54),
	.ZN(n1371));
   NAND2_X1 U1915 (.A1(REGISTERS[264]),
	.A2(n4036),
	.ZN(n351));
   OAI21_X1 U1916 (.A(n352),
	.B1(n4036),
	.B2(n56),
	.ZN(n1372));
   NAND2_X1 U1917 (.A1(REGISTERS[265]),
	.A2(n4036),
	.ZN(n352));
   OAI21_X1 U1918 (.A(n353),
	.B1(n4036),
	.B2(n58),
	.ZN(n1373));
   NAND2_X1 U1919 (.A1(REGISTERS[266]),
	.A2(n4036),
	.ZN(n353));
   OAI21_X1 U1920 (.A(n354),
	.B1(n4036),
	.B2(n60),
	.ZN(n1374));
   NAND2_X1 U1921 (.A1(REGISTERS[267]),
	.A2(FE_OFN60_n4036),
	.ZN(n354));
   OAI21_X1 U1922 (.A(n355),
	.B1(n4036),
	.B2(n62),
	.ZN(n1375));
   NAND2_X1 U1923 (.A1(REGISTERS[268]),
	.A2(n4036),
	.ZN(n355));
   OAI21_X1 U1924 (.A(n357),
	.B1(FE_OFN60_n4036),
	.B2(n66),
	.ZN(n1377));
   NAND2_X1 U1925 (.A1(REGISTERS[270]),
	.A2(FE_OFN60_n4036),
	.ZN(n357));
   OAI21_X1 U1926 (.A(n358),
	.B1(n4036),
	.B2(n68),
	.ZN(n1378));
   NAND2_X1 U1927 (.A1(REGISTERS[271]),
	.A2(n4036),
	.ZN(n358));
   OAI21_X1 U1928 (.A(n384),
	.B1(FE_OFN80_n4035),
	.B2(n52),
	.ZN(n1402));
   NAND2_X1 U1929 (.A1(REGISTERS[295]),
	.A2(FE_OFN80_n4035),
	.ZN(n384));
   OAI21_X1 U1930 (.A(n385),
	.B1(n4035),
	.B2(n54),
	.ZN(n1403));
   NAND2_X1 U1931 (.A1(REGISTERS[296]),
	.A2(n4035),
	.ZN(n385));
   OAI21_X1 U1932 (.A(n386),
	.B1(FE_OFN80_n4035),
	.B2(n56),
	.ZN(n1404));
   NAND2_X1 U1933 (.A1(REGISTERS[297]),
	.A2(FE_OFN80_n4035),
	.ZN(n386));
   OAI21_X1 U1934 (.A(n387),
	.B1(n4035),
	.B2(n58),
	.ZN(n1405));
   NAND2_X1 U1935 (.A1(REGISTERS[298]),
	.A2(n4035),
	.ZN(n387));
   OAI21_X1 U1936 (.A(n388),
	.B1(FE_OFN80_n4035),
	.B2(n60),
	.ZN(n1406));
   NAND2_X1 U1937 (.A1(REGISTERS[299]),
	.A2(FE_OFN80_n4035),
	.ZN(n388));
   OAI21_X1 U1938 (.A(n389),
	.B1(n4035),
	.B2(n62),
	.ZN(n1407));
   NAND2_X1 U1939 (.A1(REGISTERS[300]),
	.A2(n4035),
	.ZN(n389));
   OAI21_X1 U1940 (.A(n391),
	.B1(FE_OFN80_n4035),
	.B2(n66),
	.ZN(n1409));
   NAND2_X1 U1941 (.A1(REGISTERS[302]),
	.A2(FE_OFN80_n4035),
	.ZN(n391));
   OAI21_X1 U1942 (.A(n392),
	.B1(n4035),
	.B2(n68),
	.ZN(n1410));
   NAND2_X1 U1943 (.A1(REGISTERS[303]),
	.A2(n4035),
	.ZN(n392));
   OAI21_X1 U1944 (.A(n417),
	.B1(FE_OFN59_n4034),
	.B2(n52),
	.ZN(n1434));
   NAND2_X1 U1945 (.A1(REGISTERS[327]),
	.A2(FE_OFN59_n4034),
	.ZN(n417));
   OAI21_X1 U1946 (.A(n418),
	.B1(FE_OFN59_n4034),
	.B2(n54),
	.ZN(n1435));
   NAND2_X1 U1947 (.A1(REGISTERS[328]),
	.A2(FE_OFN59_n4034),
	.ZN(n418));
   OAI21_X1 U1948 (.A(n419),
	.B1(n4034),
	.B2(n56),
	.ZN(n1436));
   NAND2_X1 U1949 (.A1(REGISTERS[329]),
	.A2(n4034),
	.ZN(n419));
   OAI21_X1 U1950 (.A(n420),
	.B1(FE_OFN59_n4034),
	.B2(n58),
	.ZN(n1437));
   NAND2_X1 U1951 (.A1(REGISTERS[330]),
	.A2(FE_OFN59_n4034),
	.ZN(n420));
   OAI21_X1 U1952 (.A(n421),
	.B1(n4034),
	.B2(n60),
	.ZN(n1438));
   NAND2_X1 U1953 (.A1(REGISTERS[331]),
	.A2(n4034),
	.ZN(n421));
   OAI21_X1 U1954 (.A(n422),
	.B1(FE_OFN59_n4034),
	.B2(n62),
	.ZN(n1439));
   NAND2_X1 U1955 (.A1(REGISTERS[332]),
	.A2(FE_OFN59_n4034),
	.ZN(n422));
   OAI21_X1 U1956 (.A(n424),
	.B1(n4034),
	.B2(n66),
	.ZN(n1441));
   NAND2_X1 U1957 (.A1(REGISTERS[334]),
	.A2(n4034),
	.ZN(n424));
   OAI21_X1 U1958 (.A(n425),
	.B1(n4034),
	.B2(n68),
	.ZN(n1442));
   NAND2_X1 U1959 (.A1(REGISTERS[335]),
	.A2(n4034),
	.ZN(n425));
   OAI21_X1 U1960 (.A(n450),
	.B1(FE_OFN70_n4033),
	.B2(n52),
	.ZN(n1466));
   NAND2_X1 U1961 (.A1(REGISTERS[359]),
	.A2(FE_OFN70_n4033),
	.ZN(n450));
   OAI21_X1 U1962 (.A(n451),
	.B1(FE_OFN70_n4033),
	.B2(n54),
	.ZN(n1467));
   NAND2_X1 U1963 (.A1(REGISTERS[360]),
	.A2(FE_OFN70_n4033),
	.ZN(n451));
   OAI21_X1 U1964 (.A(n452),
	.B1(n4033),
	.B2(n56),
	.ZN(n1468));
   NAND2_X1 U1965 (.A1(REGISTERS[361]),
	.A2(n4033),
	.ZN(n452));
   OAI21_X1 U1966 (.A(n453),
	.B1(FE_OFN70_n4033),
	.B2(n58),
	.ZN(n1469));
   NAND2_X1 U1967 (.A1(REGISTERS[362]),
	.A2(FE_OFN70_n4033),
	.ZN(n453));
   OAI21_X1 U1968 (.A(n454),
	.B1(n4033),
	.B2(n60),
	.ZN(n1470));
   NAND2_X1 U1969 (.A1(REGISTERS[363]),
	.A2(n4033),
	.ZN(n454));
   OAI21_X1 U1970 (.A(n455),
	.B1(FE_OFN70_n4033),
	.B2(n62),
	.ZN(n1471));
   NAND2_X1 U1971 (.A1(REGISTERS[364]),
	.A2(FE_OFN70_n4033),
	.ZN(n455));
   OAI21_X1 U1972 (.A(n457),
	.B1(n4033),
	.B2(n66),
	.ZN(n1473));
   NAND2_X1 U1973 (.A1(REGISTERS[366]),
	.A2(n4033),
	.ZN(n457));
   OAI21_X1 U1974 (.A(n458),
	.B1(n4033),
	.B2(n68),
	.ZN(n1474));
   NAND2_X1 U1975 (.A1(REGISTERS[367]),
	.A2(n4033),
	.ZN(n458));
   OAI21_X1 U1976 (.A(n483),
	.B1(FE_OFN87_n4032),
	.B2(n52),
	.ZN(n1498));
   NAND2_X1 U1977 (.A1(REGISTERS[391]),
	.A2(FE_OFN87_n4032),
	.ZN(n483));
   OAI21_X1 U1978 (.A(n484),
	.B1(n4032),
	.B2(n54),
	.ZN(n1499));
   NAND2_X1 U1979 (.A1(REGISTERS[392]),
	.A2(n4032),
	.ZN(n484));
   OAI21_X1 U1980 (.A(n485),
	.B1(FE_OFN87_n4032),
	.B2(n56),
	.ZN(n1500));
   NAND2_X1 U1981 (.A1(REGISTERS[393]),
	.A2(FE_OFN87_n4032),
	.ZN(n485));
   OAI21_X1 U1982 (.A(n486),
	.B1(n4032),
	.B2(n58),
	.ZN(n1501));
   NAND2_X1 U1983 (.A1(REGISTERS[394]),
	.A2(n4032),
	.ZN(n486));
   OAI21_X1 U1984 (.A(n487),
	.B1(FE_OFN87_n4032),
	.B2(n60),
	.ZN(n1502));
   NAND2_X1 U1985 (.A1(REGISTERS[395]),
	.A2(FE_OFN87_n4032),
	.ZN(n487));
   OAI21_X1 U1986 (.A(n488),
	.B1(n4032),
	.B2(n62),
	.ZN(n1503));
   NAND2_X1 U1987 (.A1(REGISTERS[396]),
	.A2(n4032),
	.ZN(n488));
   OAI21_X1 U1988 (.A(n490),
	.B1(FE_OFN87_n4032),
	.B2(n66),
	.ZN(n1505));
   NAND2_X1 U1989 (.A1(REGISTERS[398]),
	.A2(FE_OFN87_n4032),
	.ZN(n490));
   OAI21_X1 U1990 (.A(n491),
	.B1(n4032),
	.B2(n68),
	.ZN(n1506));
   NAND2_X1 U1991 (.A1(REGISTERS[399]),
	.A2(n4032),
	.ZN(n491));
   OAI21_X1 U1992 (.A(n516),
	.B1(FE_OFN63_n4031),
	.B2(n52),
	.ZN(n1530));
   NAND2_X1 U1993 (.A1(REGISTERS[423]),
	.A2(FE_OFN63_n4031),
	.ZN(n516));
   OAI21_X1 U1994 (.A(n517),
	.B1(FE_OFN63_n4031),
	.B2(n54),
	.ZN(n1531));
   NAND2_X1 U1995 (.A1(REGISTERS[424]),
	.A2(FE_OFN63_n4031),
	.ZN(n517));
   OAI21_X1 U1996 (.A(n518),
	.B1(n4031),
	.B2(n56),
	.ZN(n1532));
   NAND2_X1 U1997 (.A1(REGISTERS[425]),
	.A2(n4031),
	.ZN(n518));
   OAI21_X1 U1998 (.A(n519),
	.B1(FE_OFN63_n4031),
	.B2(n58),
	.ZN(n1533));
   NAND2_X1 U1999 (.A1(REGISTERS[426]),
	.A2(FE_OFN63_n4031),
	.ZN(n519));
   OAI21_X1 U2000 (.A(n520),
	.B1(n4031),
	.B2(n60),
	.ZN(n1534));
   NAND2_X1 U2001 (.A1(REGISTERS[427]),
	.A2(n4031),
	.ZN(n520));
   OAI21_X1 U2002 (.A(n521),
	.B1(FE_OFN63_n4031),
	.B2(n62),
	.ZN(n1535));
   NAND2_X1 U2003 (.A1(REGISTERS[428]),
	.A2(FE_OFN63_n4031),
	.ZN(n521));
   OAI21_X1 U2004 (.A(n523),
	.B1(FE_OFN63_n4031),
	.B2(n66),
	.ZN(n1537));
   NAND2_X1 U2005 (.A1(REGISTERS[430]),
	.A2(FE_OFN63_n4031),
	.ZN(n523));
   OAI21_X1 U2006 (.A(n524),
	.B1(n4031),
	.B2(n68),
	.ZN(n1538));
   NAND2_X1 U2007 (.A1(REGISTERS[431]),
	.A2(n4031),
	.ZN(n524));
   OAI21_X1 U2008 (.A(n549),
	.B1(FE_OFN81_n4030),
	.B2(n52),
	.ZN(n1562));
   NAND2_X1 U2009 (.A1(REGISTERS[455]),
	.A2(FE_OFN81_n4030),
	.ZN(n549));
   OAI21_X1 U2010 (.A(n550),
	.B1(n4030),
	.B2(n54),
	.ZN(n1563));
   NAND2_X1 U2011 (.A1(REGISTERS[456]),
	.A2(n4030),
	.ZN(n550));
   OAI21_X1 U2012 (.A(n551),
	.B1(FE_OFN81_n4030),
	.B2(n56),
	.ZN(n1564));
   NAND2_X1 U2013 (.A1(REGISTERS[457]),
	.A2(FE_OFN81_n4030),
	.ZN(n551));
   OAI21_X1 U2014 (.A(n552),
	.B1(n4030),
	.B2(n58),
	.ZN(n1565));
   NAND2_X1 U2015 (.A1(REGISTERS[458]),
	.A2(n4030),
	.ZN(n552));
   OAI21_X1 U2016 (.A(n553),
	.B1(FE_OFN81_n4030),
	.B2(n60),
	.ZN(n1566));
   NAND2_X1 U2017 (.A1(REGISTERS[459]),
	.A2(FE_OFN81_n4030),
	.ZN(n553));
   OAI21_X1 U2018 (.A(n554),
	.B1(n4030),
	.B2(n62),
	.ZN(n1567));
   NAND2_X1 U2019 (.A1(REGISTERS[460]),
	.A2(n4030),
	.ZN(n554));
   OAI21_X1 U2020 (.A(n556),
	.B1(FE_OFN81_n4030),
	.B2(n66),
	.ZN(n1569));
   NAND2_X1 U2021 (.A1(REGISTERS[462]),
	.A2(FE_OFN81_n4030),
	.ZN(n556));
   OAI21_X1 U2022 (.A(n557),
	.B1(n4030),
	.B2(n68),
	.ZN(n1570));
   NAND2_X1 U2023 (.A1(REGISTERS[463]),
	.A2(n4030),
	.ZN(n557));
   OAI21_X1 U2024 (.A(n582),
	.B1(FE_OFN67_n4029),
	.B2(n52),
	.ZN(n1594));
   NAND2_X1 U2025 (.A1(REGISTERS[487]),
	.A2(FE_OFN67_n4029),
	.ZN(n582));
   OAI21_X1 U2026 (.A(n583),
	.B1(n4029),
	.B2(n54),
	.ZN(n1595));
   NAND2_X1 U2027 (.A1(REGISTERS[488]),
	.A2(n4029),
	.ZN(n583));
   OAI21_X1 U2028 (.A(n584),
	.B1(FE_OFN67_n4029),
	.B2(n56),
	.ZN(n1596));
   NAND2_X1 U2029 (.A1(REGISTERS[489]),
	.A2(FE_OFN67_n4029),
	.ZN(n584));
   OAI21_X1 U2030 (.A(n585),
	.B1(n4029),
	.B2(n58),
	.ZN(n1597));
   NAND2_X1 U2031 (.A1(REGISTERS[490]),
	.A2(n4029),
	.ZN(n585));
   OAI21_X1 U2032 (.A(n586),
	.B1(FE_OFN67_n4029),
	.B2(n60),
	.ZN(n1598));
   NAND2_X1 U2033 (.A1(REGISTERS[491]),
	.A2(FE_OFN67_n4029),
	.ZN(n586));
   OAI21_X1 U2034 (.A(n587),
	.B1(n4029),
	.B2(n62),
	.ZN(n1599));
   NAND2_X1 U2035 (.A1(REGISTERS[492]),
	.A2(n4029),
	.ZN(n587));
   OAI21_X1 U2036 (.A(n589),
	.B1(FE_OFN67_n4029),
	.B2(n66),
	.ZN(n1601));
   NAND2_X1 U2037 (.A1(REGISTERS[494]),
	.A2(FE_OFN67_n4029),
	.ZN(n589));
   OAI21_X1 U2038 (.A(n590),
	.B1(n4029),
	.B2(n68),
	.ZN(n1602));
   NAND2_X1 U2039 (.A1(REGISTERS[495]),
	.A2(n4029),
	.ZN(n590));
   OAI21_X1 U2040 (.A(n615),
	.B1(FE_OFN61_n4019),
	.B2(n52),
	.ZN(n1626));
   NAND2_X1 U2041 (.A1(REGISTERS[519]),
	.A2(FE_OFN61_n4019),
	.ZN(n615));
   OAI21_X1 U2042 (.A(n616),
	.B1(n4019),
	.B2(n54),
	.ZN(n1627));
   NAND2_X1 U2043 (.A1(REGISTERS[520]),
	.A2(n4019),
	.ZN(n616));
   OAI21_X1 U2044 (.A(n617),
	.B1(n4019),
	.B2(n56),
	.ZN(n1628));
   NAND2_X1 U2045 (.A1(REGISTERS[521]),
	.A2(n4019),
	.ZN(n617));
   OAI21_X1 U2046 (.A(n618),
	.B1(n4019),
	.B2(n58),
	.ZN(n1629));
   NAND2_X1 U2047 (.A1(REGISTERS[522]),
	.A2(n4019),
	.ZN(n618));
   OAI21_X1 U2048 (.A(n619),
	.B1(n4019),
	.B2(n60),
	.ZN(n1630));
   NAND2_X1 U2049 (.A1(REGISTERS[523]),
	.A2(n4019),
	.ZN(n619));
   OAI21_X1 U2050 (.A(n620),
	.B1(n4019),
	.B2(n62),
	.ZN(n1631));
   NAND2_X1 U2051 (.A1(REGISTERS[524]),
	.A2(n4019),
	.ZN(n620));
   OAI21_X1 U2052 (.A(n622),
	.B1(FE_OFN61_n4019),
	.B2(n66),
	.ZN(n1633));
   NAND2_X1 U2053 (.A1(REGISTERS[526]),
	.A2(FE_OFN61_n4019),
	.ZN(n622));
   OAI21_X1 U2054 (.A(n623),
	.B1(FE_OFN61_n4019),
	.B2(n68),
	.ZN(n1634));
   NAND2_X1 U2055 (.A1(REGISTERS[527]),
	.A2(FE_OFN61_n4019),
	.ZN(n623));
   OAI21_X1 U2056 (.A(n649),
	.B1(FE_OFN65_n4018),
	.B2(n52),
	.ZN(n1658));
   NAND2_X1 U2057 (.A1(REGISTERS[551]),
	.A2(FE_OFN65_n4018),
	.ZN(n649));
   OAI21_X1 U2058 (.A(n650),
	.B1(FE_OFN65_n4018),
	.B2(n54),
	.ZN(n1659));
   NAND2_X1 U2059 (.A1(REGISTERS[552]),
	.A2(FE_OFN65_n4018),
	.ZN(n650));
   OAI21_X1 U2060 (.A(n651),
	.B1(n4018),
	.B2(n56),
	.ZN(n1660));
   NAND2_X1 U2061 (.A1(REGISTERS[553]),
	.A2(n4018),
	.ZN(n651));
   OAI21_X1 U2062 (.A(n652),
	.B1(FE_OFN65_n4018),
	.B2(n58),
	.ZN(n1661));
   NAND2_X1 U2063 (.A1(REGISTERS[554]),
	.A2(FE_OFN65_n4018),
	.ZN(n652));
   OAI21_X1 U2064 (.A(n653),
	.B1(n4018),
	.B2(n60),
	.ZN(n1662));
   NAND2_X1 U2065 (.A1(REGISTERS[555]),
	.A2(n4018),
	.ZN(n653));
   OAI21_X1 U2066 (.A(n654),
	.B1(FE_OFN65_n4018),
	.B2(n62),
	.ZN(n1663));
   NAND2_X1 U2067 (.A1(REGISTERS[556]),
	.A2(FE_OFN65_n4018),
	.ZN(n654));
   OAI21_X1 U2068 (.A(n656),
	.B1(FE_OFN65_n4018),
	.B2(n66),
	.ZN(n1665));
   NAND2_X1 U2069 (.A1(REGISTERS[558]),
	.A2(FE_OFN65_n4018),
	.ZN(n656));
   OAI21_X1 U2070 (.A(n657),
	.B1(n4018),
	.B2(n68),
	.ZN(n1666));
   NAND2_X1 U2071 (.A1(REGISTERS[559]),
	.A2(n4018),
	.ZN(n657));
   OAI21_X1 U2072 (.A(n682),
	.B1(FE_OFN66_n4017),
	.B2(n52),
	.ZN(n1690));
   NAND2_X1 U2073 (.A1(REGISTERS[583]),
	.A2(FE_OFN66_n4017),
	.ZN(n682));
   OAI21_X1 U2074 (.A(n683),
	.B1(n4017),
	.B2(n54),
	.ZN(n1691));
   NAND2_X1 U2075 (.A1(REGISTERS[584]),
	.A2(n4017),
	.ZN(n683));
   OAI21_X1 U2076 (.A(n684),
	.B1(FE_OFN66_n4017),
	.B2(n56),
	.ZN(n1692));
   NAND2_X1 U2077 (.A1(REGISTERS[585]),
	.A2(FE_OFN66_n4017),
	.ZN(n684));
   OAI21_X1 U2078 (.A(n685),
	.B1(n4017),
	.B2(n58),
	.ZN(n1693));
   NAND2_X1 U2079 (.A1(REGISTERS[586]),
	.A2(n4017),
	.ZN(n685));
   OAI21_X1 U2080 (.A(n686),
	.B1(FE_OFN66_n4017),
	.B2(n60),
	.ZN(n1694));
   NAND2_X1 U2081 (.A1(REGISTERS[587]),
	.A2(FE_OFN66_n4017),
	.ZN(n686));
   OAI21_X1 U2082 (.A(n687),
	.B1(n4017),
	.B2(n62),
	.ZN(n1695));
   NAND2_X1 U2083 (.A1(REGISTERS[588]),
	.A2(n4017),
	.ZN(n687));
   OAI21_X1 U2084 (.A(n689),
	.B1(FE_OFN66_n4017),
	.B2(n66),
	.ZN(n1697));
   NAND2_X1 U2085 (.A1(REGISTERS[590]),
	.A2(FE_OFN66_n4017),
	.ZN(n689));
   OAI21_X1 U2086 (.A(n690),
	.B1(FE_OFN66_n4017),
	.B2(n68),
	.ZN(n1698));
   NAND2_X1 U2087 (.A1(REGISTERS[591]),
	.A2(FE_OFN66_n4017),
	.ZN(n690));
   OAI21_X1 U2088 (.A(n715),
	.B1(FE_OFN62_n4016),
	.B2(n52),
	.ZN(n1722));
   NAND2_X1 U2089 (.A1(REGISTERS[615]),
	.A2(FE_OFN62_n4016),
	.ZN(n715));
   OAI21_X1 U2090 (.A(n716),
	.B1(FE_OFN62_n4016),
	.B2(n54),
	.ZN(n1723));
   NAND2_X1 U2091 (.A1(REGISTERS[616]),
	.A2(FE_OFN62_n4016),
	.ZN(n716));
   OAI21_X1 U2092 (.A(n717),
	.B1(n4016),
	.B2(n56),
	.ZN(n1724));
   NAND2_X1 U2093 (.A1(REGISTERS[617]),
	.A2(n4016),
	.ZN(n717));
   OAI21_X1 U2094 (.A(n718),
	.B1(FE_OFN62_n4016),
	.B2(n58),
	.ZN(n1725));
   NAND2_X1 U2095 (.A1(REGISTERS[618]),
	.A2(FE_OFN62_n4016),
	.ZN(n718));
   OAI21_X1 U2096 (.A(n719),
	.B1(n4016),
	.B2(n60),
	.ZN(n1726));
   NAND2_X1 U2097 (.A1(REGISTERS[619]),
	.A2(n4016),
	.ZN(n719));
   OAI21_X1 U2098 (.A(n720),
	.B1(FE_OFN62_n4016),
	.B2(n62),
	.ZN(n1727));
   NAND2_X1 U2099 (.A1(REGISTERS[620]),
	.A2(FE_OFN62_n4016),
	.ZN(n720));
   OAI21_X1 U2100 (.A(n722),
	.B1(FE_OFN62_n4016),
	.B2(n66),
	.ZN(n1729));
   NAND2_X1 U2101 (.A1(REGISTERS[622]),
	.A2(FE_OFN62_n4016),
	.ZN(n722));
   OAI21_X1 U2102 (.A(n723),
	.B1(n4016),
	.B2(n68),
	.ZN(n1730));
   NAND2_X1 U2103 (.A1(REGISTERS[623]),
	.A2(n4016),
	.ZN(n723));
   OAI21_X1 U2104 (.A(n748),
	.B1(FE_OFN74_n4015),
	.B2(n52),
	.ZN(n1754));
   NAND2_X1 U2105 (.A1(REGISTERS[647]),
	.A2(FE_OFN74_n4015),
	.ZN(n748));
   OAI21_X1 U2106 (.A(n749),
	.B1(n4015),
	.B2(n54),
	.ZN(n1755));
   NAND2_X1 U2107 (.A1(REGISTERS[648]),
	.A2(n4015),
	.ZN(n749));
   OAI21_X1 U2108 (.A(n750),
	.B1(n4015),
	.B2(n56),
	.ZN(n1756));
   NAND2_X1 U2109 (.A1(REGISTERS[649]),
	.A2(FE_OFN74_n4015),
	.ZN(n750));
   OAI21_X1 U2110 (.A(n751),
	.B1(n4015),
	.B2(n58),
	.ZN(n1757));
   NAND2_X1 U2111 (.A1(REGISTERS[650]),
	.A2(n4015),
	.ZN(n751));
   OAI21_X1 U2112 (.A(n752),
	.B1(FE_OFN74_n4015),
	.B2(n60),
	.ZN(n1758));
   NAND2_X1 U2113 (.A1(REGISTERS[651]),
	.A2(FE_OFN74_n4015),
	.ZN(n752));
   OAI21_X1 U2114 (.A(n753),
	.B1(n4015),
	.B2(n62),
	.ZN(n1759));
   NAND2_X1 U2115 (.A1(REGISTERS[652]),
	.A2(n4015),
	.ZN(n753));
   OAI21_X1 U2116 (.A(n755),
	.B1(FE_OFN74_n4015),
	.B2(n66),
	.ZN(n1761));
   NAND2_X1 U2117 (.A1(REGISTERS[654]),
	.A2(FE_OFN74_n4015),
	.ZN(n755));
   OAI21_X1 U2118 (.A(n756),
	.B1(FE_OFN74_n4015),
	.B2(n68),
	.ZN(n1762));
   NAND2_X1 U2119 (.A1(REGISTERS[655]),
	.A2(FE_OFN74_n4015),
	.ZN(n756));
   OAI21_X1 U2120 (.A(n781),
	.B1(FE_OFN78_n4014),
	.B2(n52),
	.ZN(n1786));
   NAND2_X1 U2121 (.A1(REGISTERS[679]),
	.A2(FE_OFN78_n4014),
	.ZN(n781));
   OAI21_X1 U2122 (.A(n782),
	.B1(n4014),
	.B2(n54),
	.ZN(n1787));
   NAND2_X1 U2123 (.A1(REGISTERS[680]),
	.A2(n4014),
	.ZN(n782));
   OAI21_X1 U2124 (.A(n783),
	.B1(n4014),
	.B2(n56),
	.ZN(n1788));
   NAND2_X1 U2125 (.A1(REGISTERS[681]),
	.A2(n4014),
	.ZN(n783));
   OAI21_X1 U2126 (.A(n784),
	.B1(n4014),
	.B2(n58),
	.ZN(n1789));
   NAND2_X1 U2127 (.A1(REGISTERS[682]),
	.A2(n4014),
	.ZN(n784));
   OAI21_X1 U2128 (.A(n785),
	.B1(n4014),
	.B2(n60),
	.ZN(n1790));
   NAND2_X1 U2129 (.A1(REGISTERS[683]),
	.A2(n4014),
	.ZN(n785));
   OAI21_X1 U2130 (.A(n786),
	.B1(n4014),
	.B2(n62),
	.ZN(n1791));
   NAND2_X1 U2131 (.A1(REGISTERS[684]),
	.A2(n4014),
	.ZN(n786));
   OAI21_X1 U2132 (.A(n788),
	.B1(FE_OFN78_n4014),
	.B2(n66),
	.ZN(n1793));
   NAND2_X1 U2133 (.A1(REGISTERS[686]),
	.A2(FE_OFN78_n4014),
	.ZN(n788));
   OAI21_X1 U2134 (.A(n789),
	.B1(FE_OFN78_n4014),
	.B2(n68),
	.ZN(n1794));
   NAND2_X1 U2135 (.A1(REGISTERS[687]),
	.A2(FE_OFN78_n4014),
	.ZN(n789));
   OAI21_X1 U2136 (.A(n814),
	.B1(FE_OFN76_n4013),
	.B2(n52),
	.ZN(n1818));
   NAND2_X1 U2137 (.A1(REGISTERS[711]),
	.A2(FE_OFN76_n4013),
	.ZN(n814));
   OAI21_X1 U2138 (.A(n815),
	.B1(n4013),
	.B2(n54),
	.ZN(n1819));
   NAND2_X1 U2139 (.A1(REGISTERS[712]),
	.A2(n4013),
	.ZN(n815));
   OAI21_X1 U2140 (.A(n816),
	.B1(FE_OFN76_n4013),
	.B2(n56),
	.ZN(n1820));
   NAND2_X1 U2141 (.A1(REGISTERS[713]),
	.A2(FE_OFN76_n4013),
	.ZN(n816));
   OAI21_X1 U2142 (.A(n817),
	.B1(n4013),
	.B2(n58),
	.ZN(n1821));
   NAND2_X1 U2143 (.A1(REGISTERS[714]),
	.A2(n4013),
	.ZN(n817));
   OAI21_X1 U2144 (.A(n818),
	.B1(FE_OFN76_n4013),
	.B2(n60),
	.ZN(n1822));
   NAND2_X1 U2145 (.A1(REGISTERS[715]),
	.A2(FE_OFN76_n4013),
	.ZN(n818));
   OAI21_X1 U2146 (.A(n819),
	.B1(n4013),
	.B2(n62),
	.ZN(n1823));
   NAND2_X1 U2147 (.A1(REGISTERS[716]),
	.A2(n4013),
	.ZN(n819));
   OAI21_X1 U2148 (.A(n821),
	.B1(FE_OFN76_n4013),
	.B2(n66),
	.ZN(n1825));
   NAND2_X1 U2149 (.A1(REGISTERS[718]),
	.A2(FE_OFN76_n4013),
	.ZN(n821));
   OAI21_X1 U2150 (.A(n822),
	.B1(FE_OFN76_n4013),
	.B2(n68),
	.ZN(n1826));
   NAND2_X1 U2151 (.A1(REGISTERS[719]),
	.A2(FE_OFN76_n4013),
	.ZN(n822));
   OAI21_X1 U2152 (.A(n847),
	.B1(FE_OFN64_n4012),
	.B2(n52),
	.ZN(n1850));
   NAND2_X1 U2153 (.A1(REGISTERS[743]),
	.A2(FE_OFN64_n4012),
	.ZN(n847));
   OAI21_X1 U2154 (.A(n848),
	.B1(n4012),
	.B2(n54),
	.ZN(n1851));
   NAND2_X1 U2155 (.A1(REGISTERS[744]),
	.A2(n4012),
	.ZN(n848));
   OAI21_X1 U2156 (.A(n849),
	.B1(n4012),
	.B2(n56),
	.ZN(n1852));
   NAND2_X1 U2157 (.A1(REGISTERS[745]),
	.A2(n4012),
	.ZN(n849));
   OAI21_X1 U2158 (.A(n850),
	.B1(n4012),
	.B2(n58),
	.ZN(n1853));
   NAND2_X1 U2159 (.A1(REGISTERS[746]),
	.A2(n4012),
	.ZN(n850));
   OAI21_X1 U2160 (.A(n851),
	.B1(n4012),
	.B2(n60),
	.ZN(n1854));
   NAND2_X1 U2161 (.A1(REGISTERS[747]),
	.A2(n4012),
	.ZN(n851));
   OAI21_X1 U2162 (.A(n852),
	.B1(n4012),
	.B2(n62),
	.ZN(n1855));
   NAND2_X1 U2163 (.A1(REGISTERS[748]),
	.A2(n4012),
	.ZN(n852));
   OAI21_X1 U2164 (.A(n854),
	.B1(FE_OFN64_n4012),
	.B2(n66),
	.ZN(n1857));
   NAND2_X1 U2165 (.A1(REGISTERS[750]),
	.A2(FE_OFN64_n4012),
	.ZN(n854));
   OAI21_X1 U2166 (.A(n855),
	.B1(FE_OFN64_n4012),
	.B2(n68),
	.ZN(n1858));
   NAND2_X1 U2167 (.A1(REGISTERS[751]),
	.A2(FE_OFN64_n4012),
	.ZN(n855));
   OAI21_X1 U2168 (.A(n338),
	.B1(FE_OFN72_n4021),
	.B2(n96),
	.ZN(n1360));
   NAND2_X1 U2169 (.A1(REGISTERS[253]),
	.A2(FE_OFN72_n4021),
	.ZN(n338));
   OAI21_X1 U2170 (.A(n339),
	.B1(FE_OFN72_n4021),
	.B2(n98),
	.ZN(n1361));
   NAND2_X1 U2171 (.A1(REGISTERS[254]),
	.A2(FE_OFN72_n4021),
	.ZN(n339));
   OAI21_X1 U2172 (.A(n372),
	.B1(FE_OFN60_n4036),
	.B2(n96),
	.ZN(n1392));
   NAND2_X1 U2173 (.A1(REGISTERS[285]),
	.A2(FE_OFN60_n4036),
	.ZN(n372));
   OAI21_X1 U2174 (.A(n373),
	.B1(FE_OFN60_n4036),
	.B2(n98),
	.ZN(n1393));
   NAND2_X1 U2175 (.A1(REGISTERS[286]),
	.A2(FE_OFN60_n4036),
	.ZN(n373));
   OAI21_X1 U2176 (.A(n902),
	.B1(n4011),
	.B2(n96),
	.ZN(n1904));
   NAND2_X1 U2177 (.A1(REGISTERS[797]),
	.A2(n4011),
	.ZN(n902));
   OAI21_X1 U2178 (.A(n903),
	.B1(FE_OFN68_n4011),
	.B2(n98),
	.ZN(n1905));
   NAND2_X1 U2179 (.A1(REGISTERS[798]),
	.A2(FE_OFN68_n4011),
	.ZN(n903));
   OAI21_X1 U2180 (.A(n936),
	.B1(n4010),
	.B2(n96),
	.ZN(n1936));
   NAND2_X1 U2181 (.A1(REGISTERS[829]),
	.A2(n4010),
	.ZN(n936));
   OAI21_X1 U2182 (.A(n937),
	.B1(FE_OFN88_n4010),
	.B2(n98),
	.ZN(n1937));
   NAND2_X1 U2183 (.A1(REGISTERS[830]),
	.A2(FE_OFN88_n4010),
	.ZN(n937));
   OAI21_X1 U2184 (.A(n969),
	.B1(n4009),
	.B2(n96),
	.ZN(n1968));
   NAND2_X1 U2197 (.A1(REGISTERS[861]),
	.A2(n4009),
	.ZN(n969));
   OAI21_X1 U2198 (.A(n970),
	.B1(FE_OFN73_n4009),
	.B2(n98),
	.ZN(n1969));
   NAND2_X1 U2199 (.A1(REGISTERS[862]),
	.A2(FE_OFN73_n4009),
	.ZN(n970));
   OAI21_X1 U2200 (.A(n1002),
	.B1(n4008),
	.B2(n96),
	.ZN(n2000));
   NAND2_X1 U2201 (.A1(REGISTERS[893]),
	.A2(n4008),
	.ZN(n1002));
   OAI21_X1 U2202 (.A(n1003),
	.B1(FE_OFN86_n4008),
	.B2(n98),
	.ZN(n2001));
   NAND2_X1 U2203 (.A1(REGISTERS[894]),
	.A2(FE_OFN86_n4008),
	.ZN(n1003));
   OAI21_X1 U2204 (.A(n1035),
	.B1(n4007),
	.B2(n96),
	.ZN(n2032));
   NAND2_X1 U2205 (.A1(REGISTERS[925]),
	.A2(n4007),
	.ZN(n1035));
   OAI21_X1 U2206 (.A(n1036),
	.B1(FE_OFN82_n4007),
	.B2(n98),
	.ZN(n2033));
   NAND2_X1 U2207 (.A1(REGISTERS[926]),
	.A2(FE_OFN82_n4007),
	.ZN(n1036));
   OAI21_X1 U2208 (.A(n1068),
	.B1(FE_OFN71_n4006),
	.B2(n96),
	.ZN(n2064));
   NAND2_X1 U2209 (.A1(REGISTERS[957]),
	.A2(FE_OFN71_n4006),
	.ZN(n1068));
   OAI21_X1 U2210 (.A(n1069),
	.B1(FE_OFN71_n4006),
	.B2(n98),
	.ZN(n2065));
   NAND2_X1 U2211 (.A1(REGISTERS[958]),
	.A2(FE_OFN71_n4006),
	.ZN(n1069));
   OAI21_X1 U2212 (.A(n1101),
	.B1(n4005),
	.B2(n96),
	.ZN(n2096));
   NAND2_X1 U2213 (.A1(REGISTERS[989]),
	.A2(n4005),
	.ZN(n1101));
   OAI21_X1 U2214 (.A(n1102),
	.B1(FE_OFN84_n4005),
	.B2(n98),
	.ZN(n2097));
   NAND2_X1 U2215 (.A1(REGISTERS[990]),
	.A2(FE_OFN84_n4005),
	.ZN(n1102));
   OAI21_X1 U2216 (.A(n39),
	.B1(FE_OFN75_n4028),
	.B2(n38),
	.ZN(n1107));
   NAND2_X1 U2217 (.A1(REGISTERS[0]),
	.A2(FE_OFN75_n4028),
	.ZN(n39));
   OAI21_X1 U2218 (.A(n41),
	.B1(n4028),
	.B2(n40),
	.ZN(n1108));
   NAND2_X1 U2219 (.A1(REGISTERS[1]),
	.A2(n4028),
	.ZN(n41));
   OAI21_X1 U2220 (.A(n43),
	.B1(FE_OFN75_n4028),
	.B2(n42),
	.ZN(n1109));
   NAND2_X1 U2221 (.A1(REGISTERS[2]),
	.A2(FE_OFN75_n4028),
	.ZN(n43));
   OAI21_X1 U2222 (.A(n45),
	.B1(FE_OFN75_n4028),
	.B2(n44),
	.ZN(n1110));
   NAND2_X1 U2223 (.A1(REGISTERS[3]),
	.A2(FE_OFN75_n4028),
	.ZN(n45));
   OAI21_X1 U2224 (.A(n47),
	.B1(n4028),
	.B2(n46),
	.ZN(n1111));
   NAND2_X1 U2225 (.A1(REGISTERS[4]),
	.A2(n4028),
	.ZN(n47));
   OAI21_X1 U2226 (.A(n49),
	.B1(FE_OFN75_n4028),
	.B2(n48),
	.ZN(n1112));
   NAND2_X1 U2227 (.A1(REGISTERS[5]),
	.A2(FE_OFN75_n4028),
	.ZN(n49));
   OAI21_X1 U2228 (.A(n51),
	.B1(n4028),
	.B2(n50),
	.ZN(n1113));
   NAND2_X1 U2229 (.A1(REGISTERS[6]),
	.A2(n4028),
	.ZN(n51));
   OAI21_X1 U2230 (.A(n65),
	.B1(n4028),
	.B2(n64),
	.ZN(n1120));
   NAND2_X1 U2231 (.A1(REGISTERS[13]),
	.A2(n4028),
	.ZN(n65));
   OAI21_X1 U2232 (.A(n71),
	.B1(FE_OFN75_n4028),
	.B2(n70),
	.ZN(n1123));
   NAND2_X1 U2233 (.A1(REGISTERS[16]),
	.A2(FE_OFN75_n4028),
	.ZN(n71));
   OAI21_X1 U2234 (.A(n73),
	.B1(FE_OFN75_n4028),
	.B2(n72),
	.ZN(n1124));
   NAND2_X1 U2235 (.A1(REGISTERS[17]),
	.A2(FE_OFN75_n4028),
	.ZN(n73));
   OAI21_X1 U2236 (.A(n75),
	.B1(n4028),
	.B2(n74),
	.ZN(n1125));
   NAND2_X1 U2237 (.A1(REGISTERS[18]),
	.A2(n4028),
	.ZN(n75));
   OAI21_X1 U2238 (.A(n77),
	.B1(FE_OFN75_n4028),
	.B2(n76),
	.ZN(n1126));
   NAND2_X1 U2239 (.A1(REGISTERS[19]),
	.A2(FE_OFN75_n4028),
	.ZN(n77));
   OAI21_X1 U2240 (.A(n79),
	.B1(n4028),
	.B2(n78),
	.ZN(n1127));
   NAND2_X1 U2241 (.A1(REGISTERS[20]),
	.A2(n4028),
	.ZN(n79));
   OAI21_X1 U2242 (.A(n81),
	.B1(FE_OFN75_n4028),
	.B2(n80),
	.ZN(n1128));
   NAND2_X1 U2243 (.A1(REGISTERS[21]),
	.A2(FE_OFN75_n4028),
	.ZN(n81));
   OAI21_X1 U2244 (.A(n83),
	.B1(FE_OFN75_n4028),
	.B2(n82),
	.ZN(n1129));
   NAND2_X1 U2245 (.A1(REGISTERS[22]),
	.A2(FE_OFN75_n4028),
	.ZN(n83));
   OAI21_X1 U2246 (.A(n85),
	.B1(FE_OFN75_n4028),
	.B2(n84),
	.ZN(n1130));
   NAND2_X1 U2247 (.A1(REGISTERS[23]),
	.A2(FE_OFN75_n4028),
	.ZN(n85));
   OAI21_X1 U2248 (.A(n87),
	.B1(n4028),
	.B2(n86),
	.ZN(n1131));
   NAND2_X1 U2249 (.A1(REGISTERS[24]),
	.A2(n4028),
	.ZN(n87));
   OAI21_X1 U2250 (.A(n89),
	.B1(FE_OFN75_n4028),
	.B2(n88),
	.ZN(n1132));
   NAND2_X1 U2251 (.A1(REGISTERS[25]),
	.A2(FE_OFN75_n4028),
	.ZN(n89));
   OAI21_X1 U2252 (.A(n91),
	.B1(n4028),
	.B2(n90),
	.ZN(n1133));
   NAND2_X1 U2253 (.A1(REGISTERS[26]),
	.A2(n4028),
	.ZN(n91));
   OAI21_X1 U2254 (.A(n93),
	.B1(FE_OFN75_n4028),
	.B2(n92),
	.ZN(n1134));
   NAND2_X1 U2255 (.A1(REGISTERS[27]),
	.A2(FE_OFN75_n4028),
	.ZN(n93));
   OAI21_X1 U2256 (.A(n95),
	.B1(FE_OFN75_n4028),
	.B2(n94),
	.ZN(n1135));
   NAND2_X1 U2257 (.A1(REGISTERS[28]),
	.A2(FE_OFN75_n4028),
	.ZN(n95));
   OAI21_X1 U2258 (.A(n97),
	.B1(FE_OFN75_n4028),
	.B2(n96),
	.ZN(n1136));
   NAND2_X1 U2259 (.A1(REGISTERS[29]),
	.A2(FE_OFN75_n4028),
	.ZN(n97));
   OAI21_X1 U2260 (.A(n99),
	.B1(FE_OFN75_n4028),
	.B2(n98),
	.ZN(n1137));
   NAND2_X1 U2261 (.A1(REGISTERS[30]),
	.A2(FE_OFN75_n4028),
	.ZN(n99));
   OAI21_X1 U2262 (.A(n101),
	.B1(n4028),
	.B2(n100),
	.ZN(n1138));
   NAND2_X1 U2263 (.A1(REGISTERS[31]),
	.A2(n4028),
	.ZN(n101));
   OAI21_X1 U2264 (.A(n105),
	.B1(FE_OFN89_n4027),
	.B2(n38),
	.ZN(n1139));
   NAND2_X1 U2265 (.A1(REGISTERS[32]),
	.A2(FE_OFN89_n4027),
	.ZN(n105));
   OAI21_X1 U2266 (.A(n106),
	.B1(n4027),
	.B2(n40),
	.ZN(n1140));
   NAND2_X1 U2267 (.A1(REGISTERS[33]),
	.A2(n4027),
	.ZN(n106));
   OAI21_X1 U2268 (.A(n107),
	.B1(FE_OFN89_n4027),
	.B2(n42),
	.ZN(n1141));
   NAND2_X1 U2269 (.A1(REGISTERS[34]),
	.A2(FE_OFN89_n4027),
	.ZN(n107));
   OAI21_X1 U2270 (.A(n108),
	.B1(FE_OFN89_n4027),
	.B2(n44),
	.ZN(n1142));
   NAND2_X1 U2271 (.A1(REGISTERS[35]),
	.A2(FE_OFN89_n4027),
	.ZN(n108));
   OAI21_X1 U2272 (.A(n109),
	.B1(n4027),
	.B2(n46),
	.ZN(n1143));
   NAND2_X1 U2273 (.A1(REGISTERS[36]),
	.A2(n4027),
	.ZN(n109));
   OAI21_X1 U2274 (.A(n110),
	.B1(FE_OFN89_n4027),
	.B2(n48),
	.ZN(n1144));
   NAND2_X1 U2275 (.A1(REGISTERS[37]),
	.A2(FE_OFN89_n4027),
	.ZN(n110));
   OAI21_X1 U2276 (.A(n111),
	.B1(n4027),
	.B2(n50),
	.ZN(n1145));
   NAND2_X1 U2277 (.A1(REGISTERS[38]),
	.A2(n4027),
	.ZN(n111));
   OAI21_X1 U2278 (.A(n118),
	.B1(n4027),
	.B2(n64),
	.ZN(n1152));
   NAND2_X1 U2279 (.A1(REGISTERS[45]),
	.A2(n4027),
	.ZN(n118));
   OAI21_X1 U2280 (.A(n121),
	.B1(FE_OFN89_n4027),
	.B2(n70),
	.ZN(n1155));
   NAND2_X1 U2281 (.A1(REGISTERS[48]),
	.A2(FE_OFN89_n4027),
	.ZN(n121));
   OAI21_X1 U2282 (.A(n122),
	.B1(FE_OFN89_n4027),
	.B2(n72),
	.ZN(n1156));
   NAND2_X1 U2283 (.A1(REGISTERS[49]),
	.A2(FE_OFN89_n4027),
	.ZN(n122));
   OAI21_X1 U2284 (.A(n123),
	.B1(n4027),
	.B2(n74),
	.ZN(n1157));
   NAND2_X1 U2285 (.A1(REGISTERS[50]),
	.A2(n4027),
	.ZN(n123));
   OAI21_X1 U2286 (.A(n124),
	.B1(FE_OFN89_n4027),
	.B2(n76),
	.ZN(n1158));
   NAND2_X1 U2287 (.A1(REGISTERS[51]),
	.A2(FE_OFN89_n4027),
	.ZN(n124));
   OAI21_X1 U2288 (.A(n125),
	.B1(n4027),
	.B2(n78),
	.ZN(n1159));
   NAND2_X1 U2289 (.A1(REGISTERS[52]),
	.A2(n4027),
	.ZN(n125));
   OAI21_X1 U2290 (.A(n126),
	.B1(FE_OFN89_n4027),
	.B2(n80),
	.ZN(n1160));
   NAND2_X1 U2291 (.A1(REGISTERS[53]),
	.A2(FE_OFN89_n4027),
	.ZN(n126));
   OAI21_X1 U2292 (.A(n127),
	.B1(FE_OFN89_n4027),
	.B2(n82),
	.ZN(n1161));
   NAND2_X1 U2293 (.A1(REGISTERS[54]),
	.A2(FE_OFN89_n4027),
	.ZN(n127));
   OAI21_X1 U2294 (.A(n128),
	.B1(FE_OFN89_n4027),
	.B2(n84),
	.ZN(n1162));
   NAND2_X1 U2295 (.A1(REGISTERS[55]),
	.A2(FE_OFN89_n4027),
	.ZN(n128));
   OAI21_X1 U2296 (.A(n129),
	.B1(n4027),
	.B2(n86),
	.ZN(n1163));
   NAND2_X1 U2297 (.A1(REGISTERS[56]),
	.A2(n4027),
	.ZN(n129));
   OAI21_X1 U2298 (.A(n130),
	.B1(FE_OFN89_n4027),
	.B2(n88),
	.ZN(n1164));
   NAND2_X1 U2299 (.A1(REGISTERS[57]),
	.A2(FE_OFN89_n4027),
	.ZN(n130));
   OAI21_X1 U2300 (.A(n131),
	.B1(n4027),
	.B2(n90),
	.ZN(n1165));
   NAND2_X1 U2301 (.A1(REGISTERS[58]),
	.A2(n4027),
	.ZN(n131));
   OAI21_X1 U2302 (.A(n132),
	.B1(FE_OFN89_n4027),
	.B2(n92),
	.ZN(n1166));
   NAND2_X1 U2303 (.A1(REGISTERS[59]),
	.A2(FE_OFN89_n4027),
	.ZN(n132));
   OAI21_X1 U2304 (.A(n133),
	.B1(FE_OFN89_n4027),
	.B2(n94),
	.ZN(n1167));
   NAND2_X1 U2305 (.A1(REGISTERS[60]),
	.A2(FE_OFN89_n4027),
	.ZN(n133));
   OAI21_X1 U2306 (.A(n134),
	.B1(FE_OFN89_n4027),
	.B2(n96),
	.ZN(n1168));
   NAND2_X1 U2307 (.A1(REGISTERS[61]),
	.A2(FE_OFN89_n4027),
	.ZN(n134));
   OAI21_X1 U2308 (.A(n135),
	.B1(FE_OFN89_n4027),
	.B2(n98),
	.ZN(n1169));
   NAND2_X1 U2309 (.A1(REGISTERS[62]),
	.A2(FE_OFN89_n4027),
	.ZN(n135));
   OAI21_X1 U2310 (.A(n136),
	.B1(n4027),
	.B2(n100),
	.ZN(n1170));
   NAND2_X1 U2311 (.A1(REGISTERS[63]),
	.A2(n4027),
	.ZN(n136));
   OAI21_X1 U2312 (.A(n139),
	.B1(FE_OFN77_n4026),
	.B2(n38),
	.ZN(n1171));
   NAND2_X1 U2313 (.A1(REGISTERS[64]),
	.A2(FE_OFN77_n4026),
	.ZN(n139));
   OAI21_X1 U2314 (.A(n140),
	.B1(n4026),
	.B2(n40),
	.ZN(n1172));
   NAND2_X1 U2315 (.A1(REGISTERS[65]),
	.A2(n4026),
	.ZN(n140));
   OAI21_X1 U2316 (.A(n141),
	.B1(FE_OFN77_n4026),
	.B2(n42),
	.ZN(n1173));
   NAND2_X1 U2317 (.A1(REGISTERS[66]),
	.A2(FE_OFN77_n4026),
	.ZN(n141));
   OAI21_X1 U2318 (.A(n142),
	.B1(FE_OFN77_n4026),
	.B2(n44),
	.ZN(n1174));
   NAND2_X1 U2319 (.A1(REGISTERS[67]),
	.A2(FE_OFN77_n4026),
	.ZN(n142));
   OAI21_X1 U2320 (.A(n143),
	.B1(n4026),
	.B2(n46),
	.ZN(n1175));
   NAND2_X1 U2321 (.A1(REGISTERS[68]),
	.A2(n4026),
	.ZN(n143));
   OAI21_X1 U2322 (.A(n144),
	.B1(FE_OFN77_n4026),
	.B2(n48),
	.ZN(n1176));
   NAND2_X1 U2323 (.A1(REGISTERS[69]),
	.A2(FE_OFN77_n4026),
	.ZN(n144));
   OAI21_X1 U2324 (.A(n145),
	.B1(n4026),
	.B2(n50),
	.ZN(n1177));
   NAND2_X1 U2325 (.A1(REGISTERS[70]),
	.A2(n4026),
	.ZN(n145));
   OAI21_X1 U2326 (.A(n152),
	.B1(n4026),
	.B2(n64),
	.ZN(n1184));
   NAND2_X1 U2327 (.A1(REGISTERS[77]),
	.A2(n4026),
	.ZN(n152));
   OAI21_X1 U2328 (.A(n155),
	.B1(FE_OFN77_n4026),
	.B2(n70),
	.ZN(n1187));
   NAND2_X1 U2329 (.A1(REGISTERS[80]),
	.A2(FE_OFN77_n4026),
	.ZN(n155));
   OAI21_X1 U2330 (.A(n156),
	.B1(FE_OFN77_n4026),
	.B2(n72),
	.ZN(n1188));
   NAND2_X1 U2331 (.A1(REGISTERS[81]),
	.A2(FE_OFN77_n4026),
	.ZN(n156));
   OAI21_X1 U2332 (.A(n157),
	.B1(n4026),
	.B2(n74),
	.ZN(n1189));
   NAND2_X1 U2333 (.A1(REGISTERS[82]),
	.A2(n4026),
	.ZN(n157));
   OAI21_X1 U2334 (.A(n158),
	.B1(FE_OFN77_n4026),
	.B2(n76),
	.ZN(n1190));
   NAND2_X1 U2335 (.A1(REGISTERS[83]),
	.A2(FE_OFN77_n4026),
	.ZN(n158));
   OAI21_X1 U2336 (.A(n159),
	.B1(n4026),
	.B2(n78),
	.ZN(n1191));
   NAND2_X1 U2337 (.A1(REGISTERS[84]),
	.A2(n4026),
	.ZN(n159));
   OAI21_X1 U2338 (.A(n160),
	.B1(FE_OFN77_n4026),
	.B2(n80),
	.ZN(n1192));
   NAND2_X1 U2339 (.A1(REGISTERS[85]),
	.A2(FE_OFN77_n4026),
	.ZN(n160));
   OAI21_X1 U2340 (.A(n161),
	.B1(FE_OFN77_n4026),
	.B2(n82),
	.ZN(n1193));
   NAND2_X1 U2341 (.A1(REGISTERS[86]),
	.A2(FE_OFN77_n4026),
	.ZN(n161));
   OAI21_X1 U2342 (.A(n162),
	.B1(FE_OFN77_n4026),
	.B2(n84),
	.ZN(n1194));
   NAND2_X1 U2343 (.A1(REGISTERS[87]),
	.A2(FE_OFN77_n4026),
	.ZN(n162));
   OAI21_X1 U2344 (.A(n163),
	.B1(n4026),
	.B2(n86),
	.ZN(n1195));
   NAND2_X1 U2345 (.A1(REGISTERS[88]),
	.A2(n4026),
	.ZN(n163));
   OAI21_X1 U2346 (.A(n164),
	.B1(FE_OFN77_n4026),
	.B2(n88),
	.ZN(n1196));
   NAND2_X1 U2347 (.A1(REGISTERS[89]),
	.A2(FE_OFN77_n4026),
	.ZN(n164));
   OAI21_X1 U2348 (.A(n165),
	.B1(n4026),
	.B2(n90),
	.ZN(n1197));
   NAND2_X1 U2349 (.A1(REGISTERS[90]),
	.A2(n4026),
	.ZN(n165));
   OAI21_X1 U2350 (.A(n166),
	.B1(FE_OFN77_n4026),
	.B2(n92),
	.ZN(n1198));
   NAND2_X1 U2351 (.A1(REGISTERS[91]),
	.A2(FE_OFN77_n4026),
	.ZN(n166));
   OAI21_X1 U2352 (.A(n167),
	.B1(FE_OFN77_n4026),
	.B2(n94),
	.ZN(n1199));
   NAND2_X1 U2353 (.A1(REGISTERS[92]),
	.A2(FE_OFN77_n4026),
	.ZN(n167));
   OAI21_X1 U2354 (.A(n168),
	.B1(FE_OFN77_n4026),
	.B2(n96),
	.ZN(n1200));
   NAND2_X1 U2355 (.A1(REGISTERS[93]),
	.A2(FE_OFN77_n4026),
	.ZN(n168));
   OAI21_X1 U2356 (.A(n169),
	.B1(FE_OFN77_n4026),
	.B2(n98),
	.ZN(n1201));
   NAND2_X1 U2357 (.A1(REGISTERS[94]),
	.A2(FE_OFN77_n4026),
	.ZN(n169));
   OAI21_X1 U2358 (.A(n170),
	.B1(n4026),
	.B2(n100),
	.ZN(n1202));
   NAND2_X1 U2359 (.A1(REGISTERS[95]),
	.A2(n4026),
	.ZN(n170));
   OAI21_X1 U2360 (.A(n173),
	.B1(FE_OFN69_n4025),
	.B2(n38),
	.ZN(n1203));
   NAND2_X1 U2361 (.A1(REGISTERS[96]),
	.A2(FE_OFN69_n4025),
	.ZN(n173));
   OAI21_X1 U2362 (.A(n174),
	.B1(FE_OFN69_n4025),
	.B2(n40),
	.ZN(n1204));
   NAND2_X1 U2363 (.A1(REGISTERS[97]),
	.A2(FE_OFN69_n4025),
	.ZN(n174));
   OAI21_X1 U2364 (.A(n175),
	.B1(FE_OFN69_n4025),
	.B2(n42),
	.ZN(n1205));
   NAND2_X1 U2365 (.A1(REGISTERS[98]),
	.A2(FE_OFN69_n4025),
	.ZN(n175));
   OAI21_X1 U2366 (.A(n176),
	.B1(FE_OFN69_n4025),
	.B2(n44),
	.ZN(n1206));
   NAND2_X1 U2367 (.A1(REGISTERS[99]),
	.A2(FE_OFN69_n4025),
	.ZN(n176));
   OAI21_X1 U2368 (.A(n177),
	.B1(n4025),
	.B2(n46),
	.ZN(n1207));
   NAND2_X1 U2369 (.A1(REGISTERS[100]),
	.A2(n4025),
	.ZN(n177));
   OAI21_X1 U2370 (.A(n178),
	.B1(FE_OFN69_n4025),
	.B2(n48),
	.ZN(n1208));
   NAND2_X1 U2371 (.A1(REGISTERS[101]),
	.A2(FE_OFN69_n4025),
	.ZN(n178));
   OAI21_X1 U2372 (.A(n179),
	.B1(FE_OFN69_n4025),
	.B2(n50),
	.ZN(n1209));
   NAND2_X1 U2373 (.A1(REGISTERS[102]),
	.A2(FE_OFN69_n4025),
	.ZN(n179));
   OAI21_X1 U2374 (.A(n186),
	.B1(FE_OFN69_n4025),
	.B2(n64),
	.ZN(n1216));
   NAND2_X1 U2375 (.A1(REGISTERS[109]),
	.A2(FE_OFN69_n4025),
	.ZN(n186));
   OAI21_X1 U2376 (.A(n189),
	.B1(FE_OFN69_n4025),
	.B2(n70),
	.ZN(n1219));
   NAND2_X1 U2377 (.A1(REGISTERS[112]),
	.A2(FE_OFN69_n4025),
	.ZN(n189));
   OAI21_X1 U2378 (.A(n190),
	.B1(FE_OFN69_n4025),
	.B2(n72),
	.ZN(n1220));
   NAND2_X1 U2379 (.A1(REGISTERS[113]),
	.A2(FE_OFN69_n4025),
	.ZN(n190));
   OAI21_X1 U2380 (.A(n191),
	.B1(FE_OFN69_n4025),
	.B2(n74),
	.ZN(n1221));
   NAND2_X1 U2381 (.A1(REGISTERS[114]),
	.A2(FE_OFN69_n4025),
	.ZN(n191));
   OAI21_X1 U2382 (.A(n192),
	.B1(FE_OFN69_n4025),
	.B2(n76),
	.ZN(n1222));
   NAND2_X1 U2383 (.A1(REGISTERS[115]),
	.A2(FE_OFN69_n4025),
	.ZN(n192));
   OAI21_X1 U2384 (.A(n193),
	.B1(FE_OFN69_n4025),
	.B2(n78),
	.ZN(n1223));
   NAND2_X1 U2385 (.A1(REGISTERS[116]),
	.A2(FE_OFN69_n4025),
	.ZN(n193));
   OAI21_X1 U2386 (.A(n194),
	.B1(FE_OFN69_n4025),
	.B2(n80),
	.ZN(n1224));
   NAND2_X1 U2387 (.A1(REGISTERS[117]),
	.A2(FE_OFN69_n4025),
	.ZN(n194));
   OAI21_X1 U2388 (.A(n195),
	.B1(FE_OFN69_n4025),
	.B2(n82),
	.ZN(n1225));
   NAND2_X1 U2389 (.A1(REGISTERS[118]),
	.A2(FE_OFN69_n4025),
	.ZN(n195));
   OAI21_X1 U2390 (.A(n196),
	.B1(FE_OFN69_n4025),
	.B2(n84),
	.ZN(n1226));
   NAND2_X1 U2391 (.A1(REGISTERS[119]),
	.A2(FE_OFN69_n4025),
	.ZN(n196));
   OAI21_X1 U2392 (.A(n197),
	.B1(FE_OFN69_n4025),
	.B2(n86),
	.ZN(n1227));
   NAND2_X1 U2393 (.A1(REGISTERS[120]),
	.A2(FE_OFN69_n4025),
	.ZN(n197));
   OAI21_X1 U2394 (.A(n198),
	.B1(FE_OFN69_n4025),
	.B2(n88),
	.ZN(n1228));
   NAND2_X1 U2395 (.A1(REGISTERS[121]),
	.A2(FE_OFN69_n4025),
	.ZN(n198));
   OAI21_X1 U2396 (.A(n199),
	.B1(FE_OFN69_n4025),
	.B2(n90),
	.ZN(n1229));
   NAND2_X1 U2397 (.A1(REGISTERS[122]),
	.A2(FE_OFN69_n4025),
	.ZN(n199));
   OAI21_X1 U2398 (.A(n200),
	.B1(FE_OFN69_n4025),
	.B2(n92),
	.ZN(n1230));
   NAND2_X1 U2399 (.A1(REGISTERS[123]),
	.A2(FE_OFN69_n4025),
	.ZN(n200));
   OAI21_X1 U2400 (.A(n201),
	.B1(FE_OFN69_n4025),
	.B2(n94),
	.ZN(n1231));
   NAND2_X1 U2401 (.A1(REGISTERS[124]),
	.A2(FE_OFN69_n4025),
	.ZN(n201));
   OAI21_X1 U2402 (.A(n202),
	.B1(FE_OFN69_n4025),
	.B2(n96),
	.ZN(n1232));
   NAND2_X1 U2403 (.A1(REGISTERS[125]),
	.A2(FE_OFN69_n4025),
	.ZN(n202));
   OAI21_X1 U2404 (.A(n203),
	.B1(FE_OFN69_n4025),
	.B2(n98),
	.ZN(n1233));
   NAND2_X1 U2405 (.A1(REGISTERS[126]),
	.A2(FE_OFN69_n4025),
	.ZN(n203));
   OAI21_X1 U2406 (.A(n204),
	.B1(FE_OFN69_n4025),
	.B2(n100),
	.ZN(n1234));
   NAND2_X1 U2407 (.A1(REGISTERS[127]),
	.A2(FE_OFN69_n4025),
	.ZN(n204));
   OAI21_X1 U2408 (.A(n241),
	.B1(FE_OFN79_n4023),
	.B2(n38),
	.ZN(n1267));
   NAND2_X1 U2409 (.A1(REGISTERS[160]),
	.A2(FE_OFN79_n4023),
	.ZN(n241));
   OAI21_X1 U2410 (.A(n242),
	.B1(n4023),
	.B2(n40),
	.ZN(n1268));
   NAND2_X1 U2411 (.A1(REGISTERS[161]),
	.A2(n4023),
	.ZN(n242));
   OAI21_X1 U2412 (.A(n243),
	.B1(FE_OFN79_n4023),
	.B2(n42),
	.ZN(n1269));
   NAND2_X1 U2413 (.A1(REGISTERS[162]),
	.A2(FE_OFN79_n4023),
	.ZN(n243));
   OAI21_X1 U2414 (.A(n244),
	.B1(FE_OFN79_n4023),
	.B2(n44),
	.ZN(n1270));
   NAND2_X1 U2415 (.A1(REGISTERS[163]),
	.A2(FE_OFN79_n4023),
	.ZN(n244));
   OAI21_X1 U2416 (.A(n245),
	.B1(n4023),
	.B2(n46),
	.ZN(n1271));
   NAND2_X1 U2417 (.A1(REGISTERS[164]),
	.A2(n4023),
	.ZN(n245));
   OAI21_X1 U2418 (.A(n246),
	.B1(FE_OFN79_n4023),
	.B2(n48),
	.ZN(n1272));
   NAND2_X1 U2419 (.A1(REGISTERS[165]),
	.A2(FE_OFN79_n4023),
	.ZN(n246));
   OAI21_X1 U2420 (.A(n247),
	.B1(n4023),
	.B2(n50),
	.ZN(n1273));
   NAND2_X1 U2421 (.A1(REGISTERS[166]),
	.A2(n4023),
	.ZN(n247));
   OAI21_X1 U2422 (.A(n254),
	.B1(n4023),
	.B2(n64),
	.ZN(n1280));
   NAND2_X1 U2423 (.A1(REGISTERS[173]),
	.A2(n4023),
	.ZN(n254));
   OAI21_X1 U2424 (.A(n257),
	.B1(FE_OFN79_n4023),
	.B2(n70),
	.ZN(n1283));
   NAND2_X1 U2425 (.A1(REGISTERS[176]),
	.A2(FE_OFN79_n4023),
	.ZN(n257));
   OAI21_X1 U2426 (.A(n258),
	.B1(FE_OFN79_n4023),
	.B2(n72),
	.ZN(n1284));
   NAND2_X1 U2427 (.A1(REGISTERS[177]),
	.A2(FE_OFN79_n4023),
	.ZN(n258));
   OAI21_X1 U2428 (.A(n259),
	.B1(n4023),
	.B2(n74),
	.ZN(n1285));
   NAND2_X1 U2429 (.A1(REGISTERS[178]),
	.A2(n4023),
	.ZN(n259));
   OAI21_X1 U2430 (.A(n260),
	.B1(FE_OFN79_n4023),
	.B2(n76),
	.ZN(n1286));
   NAND2_X1 U2431 (.A1(REGISTERS[179]),
	.A2(FE_OFN79_n4023),
	.ZN(n260));
   OAI21_X1 U2432 (.A(n261),
	.B1(n4023),
	.B2(n78),
	.ZN(n1287));
   NAND2_X1 U2433 (.A1(REGISTERS[180]),
	.A2(n4023),
	.ZN(n261));
   OAI21_X1 U2434 (.A(n262),
	.B1(FE_OFN79_n4023),
	.B2(n80),
	.ZN(n1288));
   NAND2_X1 U2435 (.A1(REGISTERS[181]),
	.A2(FE_OFN79_n4023),
	.ZN(n262));
   OAI21_X1 U2436 (.A(n263),
	.B1(FE_OFN79_n4023),
	.B2(n82),
	.ZN(n1289));
   NAND2_X1 U2437 (.A1(REGISTERS[182]),
	.A2(FE_OFN79_n4023),
	.ZN(n263));
   OAI21_X1 U2438 (.A(n264),
	.B1(FE_OFN79_n4023),
	.B2(n84),
	.ZN(n1290));
   NAND2_X1 U2439 (.A1(REGISTERS[183]),
	.A2(FE_OFN79_n4023),
	.ZN(n264));
   OAI21_X1 U2440 (.A(n265),
	.B1(n4023),
	.B2(n86),
	.ZN(n1291));
   NAND2_X1 U2441 (.A1(REGISTERS[184]),
	.A2(n4023),
	.ZN(n265));
   OAI21_X1 U2442 (.A(n266),
	.B1(FE_OFN79_n4023),
	.B2(n88),
	.ZN(n1292));
   NAND2_X1 U2443 (.A1(REGISTERS[185]),
	.A2(FE_OFN79_n4023),
	.ZN(n266));
   OAI21_X1 U2444 (.A(n267),
	.B1(n4023),
	.B2(n90),
	.ZN(n1293));
   NAND2_X1 U2445 (.A1(REGISTERS[186]),
	.A2(n4023),
	.ZN(n267));
   OAI21_X1 U2446 (.A(n268),
	.B1(FE_OFN79_n4023),
	.B2(n92),
	.ZN(n1294));
   NAND2_X1 U2447 (.A1(REGISTERS[187]),
	.A2(FE_OFN79_n4023),
	.ZN(n268));
   OAI21_X1 U2448 (.A(n269),
	.B1(FE_OFN79_n4023),
	.B2(n94),
	.ZN(n1295));
   NAND2_X1 U2449 (.A1(REGISTERS[188]),
	.A2(FE_OFN79_n4023),
	.ZN(n269));
   OAI21_X1 U2450 (.A(n270),
	.B1(FE_OFN79_n4023),
	.B2(n96),
	.ZN(n1296));
   NAND2_X1 U2451 (.A1(REGISTERS[189]),
	.A2(FE_OFN79_n4023),
	.ZN(n270));
   OAI21_X1 U2452 (.A(n271),
	.B1(FE_OFN79_n4023),
	.B2(n98),
	.ZN(n1297));
   NAND2_X1 U2453 (.A1(REGISTERS[190]),
	.A2(FE_OFN79_n4023),
	.ZN(n271));
   OAI21_X1 U2454 (.A(n272),
	.B1(n4023),
	.B2(n100),
	.ZN(n1298));
   NAND2_X1 U2455 (.A1(REGISTERS[191]),
	.A2(n4023),
	.ZN(n272));
   OAI21_X1 U2456 (.A(n275),
	.B1(FE_OFN85_n4022),
	.B2(n38),
	.ZN(n1299));
   NAND2_X1 U2457 (.A1(REGISTERS[192]),
	.A2(FE_OFN85_n4022),
	.ZN(n275));
   OAI21_X1 U2458 (.A(n276),
	.B1(n4022),
	.B2(n40),
	.ZN(n1300));
   NAND2_X1 U2459 (.A1(REGISTERS[193]),
	.A2(n4022),
	.ZN(n276));
   OAI21_X1 U2460 (.A(n277),
	.B1(FE_OFN85_n4022),
	.B2(n42),
	.ZN(n1301));
   NAND2_X1 U2461 (.A1(REGISTERS[194]),
	.A2(FE_OFN85_n4022),
	.ZN(n277));
   OAI21_X1 U2462 (.A(n278),
	.B1(FE_OFN85_n4022),
	.B2(n44),
	.ZN(n1302));
   NAND2_X1 U2463 (.A1(REGISTERS[195]),
	.A2(FE_OFN85_n4022),
	.ZN(n278));
   OAI21_X1 U2464 (.A(n279),
	.B1(n4022),
	.B2(n46),
	.ZN(n1303));
   NAND2_X1 U2465 (.A1(REGISTERS[196]),
	.A2(n4022),
	.ZN(n279));
   OAI21_X1 U2466 (.A(n280),
	.B1(FE_OFN85_n4022),
	.B2(n48),
	.ZN(n1304));
   NAND2_X1 U2467 (.A1(REGISTERS[197]),
	.A2(FE_OFN85_n4022),
	.ZN(n280));
   OAI21_X1 U2468 (.A(n281),
	.B1(n4022),
	.B2(n50),
	.ZN(n1305));
   NAND2_X1 U2469 (.A1(REGISTERS[198]),
	.A2(n4022),
	.ZN(n281));
   OAI21_X1 U2470 (.A(n288),
	.B1(n4022),
	.B2(n64),
	.ZN(n1312));
   NAND2_X1 U2471 (.A1(REGISTERS[205]),
	.A2(n4022),
	.ZN(n288));
   OAI21_X1 U2472 (.A(n291),
	.B1(FE_OFN85_n4022),
	.B2(n70),
	.ZN(n1315));
   NAND2_X1 U2473 (.A1(REGISTERS[208]),
	.A2(FE_OFN85_n4022),
	.ZN(n291));
   OAI21_X1 U2474 (.A(n292),
	.B1(FE_OFN85_n4022),
	.B2(n72),
	.ZN(n1316));
   NAND2_X1 U2475 (.A1(REGISTERS[209]),
	.A2(FE_OFN85_n4022),
	.ZN(n292));
   OAI21_X1 U2476 (.A(n293),
	.B1(n4022),
	.B2(n74),
	.ZN(n1317));
   NAND2_X1 U2477 (.A1(REGISTERS[210]),
	.A2(n4022),
	.ZN(n293));
   OAI21_X1 U2478 (.A(n294),
	.B1(FE_OFN85_n4022),
	.B2(n76),
	.ZN(n1318));
   NAND2_X1 U2479 (.A1(REGISTERS[211]),
	.A2(FE_OFN85_n4022),
	.ZN(n294));
   OAI21_X1 U2480 (.A(n295),
	.B1(n4022),
	.B2(n78),
	.ZN(n1319));
   NAND2_X1 U2481 (.A1(REGISTERS[212]),
	.A2(n4022),
	.ZN(n295));
   OAI21_X1 U2482 (.A(n296),
	.B1(FE_OFN85_n4022),
	.B2(n80),
	.ZN(n1320));
   NAND2_X1 U2483 (.A1(REGISTERS[213]),
	.A2(FE_OFN85_n4022),
	.ZN(n296));
   OAI21_X1 U2484 (.A(n297),
	.B1(FE_OFN85_n4022),
	.B2(n82),
	.ZN(n1321));
   NAND2_X1 U2485 (.A1(REGISTERS[214]),
	.A2(FE_OFN85_n4022),
	.ZN(n297));
   OAI21_X1 U2486 (.A(n298),
	.B1(FE_OFN85_n4022),
	.B2(n84),
	.ZN(n1322));
   NAND2_X1 U2487 (.A1(REGISTERS[215]),
	.A2(FE_OFN85_n4022),
	.ZN(n298));
   OAI21_X1 U2488 (.A(n299),
	.B1(n4022),
	.B2(n86),
	.ZN(n1323));
   NAND2_X1 U2489 (.A1(REGISTERS[216]),
	.A2(n4022),
	.ZN(n299));
   OAI21_X1 U2490 (.A(n300),
	.B1(FE_OFN85_n4022),
	.B2(n88),
	.ZN(n1324));
   NAND2_X1 U2491 (.A1(REGISTERS[217]),
	.A2(FE_OFN85_n4022),
	.ZN(n300));
   OAI21_X1 U2492 (.A(n301),
	.B1(n4022),
	.B2(n90),
	.ZN(n1325));
   NAND2_X1 U2493 (.A1(REGISTERS[218]),
	.A2(n4022),
	.ZN(n301));
   OAI21_X1 U2494 (.A(n302),
	.B1(FE_OFN85_n4022),
	.B2(n92),
	.ZN(n1326));
   NAND2_X1 U2495 (.A1(REGISTERS[219]),
	.A2(FE_OFN85_n4022),
	.ZN(n302));
   OAI21_X1 U2496 (.A(n303),
	.B1(FE_OFN85_n4022),
	.B2(n94),
	.ZN(n1327));
   NAND2_X1 U2497 (.A1(REGISTERS[220]),
	.A2(FE_OFN85_n4022),
	.ZN(n303));
   OAI21_X1 U2498 (.A(n304),
	.B1(FE_OFN85_n4022),
	.B2(n96),
	.ZN(n1328));
   NAND2_X1 U2499 (.A1(REGISTERS[221]),
	.A2(FE_OFN85_n4022),
	.ZN(n304));
   OAI21_X1 U2500 (.A(n305),
	.B1(FE_OFN85_n4022),
	.B2(n98),
	.ZN(n1329));
   NAND2_X1 U2501 (.A1(REGISTERS[222]),
	.A2(FE_OFN85_n4022),
	.ZN(n305));
   OAI21_X1 U2502 (.A(n306),
	.B1(n4022),
	.B2(n100),
	.ZN(n1330));
   NAND2_X1 U2503 (.A1(REGISTERS[223]),
	.A2(n4022),
	.ZN(n306));
   OAI21_X1 U2504 (.A(n309),
	.B1(FE_OFN72_n4021),
	.B2(n38),
	.ZN(n1331));
   NAND2_X1 U2505 (.A1(REGISTERS[224]),
	.A2(FE_OFN72_n4021),
	.ZN(n309));
   OAI21_X1 U2506 (.A(n310),
	.B1(n4021),
	.B2(n40),
	.ZN(n1332));
   NAND2_X1 U2507 (.A1(REGISTERS[225]),
	.A2(n4021),
	.ZN(n310));
   OAI21_X1 U2508 (.A(n311),
	.B1(FE_OFN72_n4021),
	.B2(n42),
	.ZN(n1333));
   NAND2_X1 U2509 (.A1(REGISTERS[226]),
	.A2(FE_OFN72_n4021),
	.ZN(n311));
   OAI21_X1 U2510 (.A(n312),
	.B1(FE_OFN72_n4021),
	.B2(n44),
	.ZN(n1334));
   NAND2_X1 U2511 (.A1(REGISTERS[227]),
	.A2(FE_OFN72_n4021),
	.ZN(n312));
   OAI21_X1 U2512 (.A(n313),
	.B1(n4021),
	.B2(n46),
	.ZN(n1335));
   NAND2_X1 U2513 (.A1(REGISTERS[228]),
	.A2(n4021),
	.ZN(n313));
   OAI21_X1 U2514 (.A(n314),
	.B1(FE_OFN72_n4021),
	.B2(n48),
	.ZN(n1336));
   NAND2_X1 U2515 (.A1(REGISTERS[229]),
	.A2(FE_OFN72_n4021),
	.ZN(n314));
   OAI21_X1 U2516 (.A(n315),
	.B1(n4021),
	.B2(n50),
	.ZN(n1337));
   NAND2_X1 U2517 (.A1(REGISTERS[230]),
	.A2(n4021),
	.ZN(n315));
   OAI21_X1 U2518 (.A(n322),
	.B1(n4021),
	.B2(n64),
	.ZN(n1344));
   NAND2_X1 U2519 (.A1(REGISTERS[237]),
	.A2(n4021),
	.ZN(n322));
   OAI21_X1 U2520 (.A(n325),
	.B1(FE_OFN72_n4021),
	.B2(n70),
	.ZN(n1347));
   NAND2_X1 U2521 (.A1(REGISTERS[240]),
	.A2(FE_OFN72_n4021),
	.ZN(n325));
   OAI21_X1 U2522 (.A(n326),
	.B1(FE_OFN72_n4021),
	.B2(n72),
	.ZN(n1348));
   NAND2_X1 U2523 (.A1(REGISTERS[241]),
	.A2(FE_OFN72_n4021),
	.ZN(n326));
   OAI21_X1 U2524 (.A(n327),
	.B1(n4021),
	.B2(n74),
	.ZN(n1349));
   NAND2_X1 U2525 (.A1(REGISTERS[242]),
	.A2(n4021),
	.ZN(n327));
   OAI21_X1 U2526 (.A(n328),
	.B1(FE_OFN72_n4021),
	.B2(n76),
	.ZN(n1350));
   NAND2_X1 U2527 (.A1(REGISTERS[243]),
	.A2(FE_OFN72_n4021),
	.ZN(n328));
   OAI21_X1 U2528 (.A(n329),
	.B1(n4021),
	.B2(n78),
	.ZN(n1351));
   NAND2_X1 U2529 (.A1(REGISTERS[244]),
	.A2(n4021),
	.ZN(n329));
   OAI21_X1 U2530 (.A(n330),
	.B1(FE_OFN72_n4021),
	.B2(n80),
	.ZN(n1352));
   NAND2_X1 U2531 (.A1(REGISTERS[245]),
	.A2(FE_OFN72_n4021),
	.ZN(n330));
   OAI21_X1 U2532 (.A(n331),
	.B1(FE_OFN72_n4021),
	.B2(n82),
	.ZN(n1353));
   NAND2_X1 U2533 (.A1(REGISTERS[246]),
	.A2(FE_OFN72_n4021),
	.ZN(n331));
   OAI21_X1 U2534 (.A(n332),
	.B1(FE_OFN72_n4021),
	.B2(n84),
	.ZN(n1354));
   NAND2_X1 U2535 (.A1(REGISTERS[247]),
	.A2(FE_OFN72_n4021),
	.ZN(n332));
   OAI21_X1 U2536 (.A(n333),
	.B1(n4021),
	.B2(n86),
	.ZN(n1355));
   NAND2_X1 U2537 (.A1(REGISTERS[248]),
	.A2(n4021),
	.ZN(n333));
   OAI21_X1 U2538 (.A(n334),
	.B1(FE_OFN72_n4021),
	.B2(n88),
	.ZN(n1356));
   NAND2_X1 U2539 (.A1(REGISTERS[249]),
	.A2(FE_OFN72_n4021),
	.ZN(n334));
   OAI21_X1 U2540 (.A(n335),
	.B1(n4021),
	.B2(n90),
	.ZN(n1357));
   NAND2_X1 U2541 (.A1(REGISTERS[250]),
	.A2(n4021),
	.ZN(n335));
   OAI21_X1 U2542 (.A(n336),
	.B1(FE_OFN72_n4021),
	.B2(n92),
	.ZN(n1358));
   NAND2_X1 U2543 (.A1(REGISTERS[251]),
	.A2(FE_OFN72_n4021),
	.ZN(n336));
   OAI21_X1 U2544 (.A(n337),
	.B1(FE_OFN72_n4021),
	.B2(n94),
	.ZN(n1359));
   NAND2_X1 U2545 (.A1(REGISTERS[252]),
	.A2(FE_OFN72_n4021),
	.ZN(n337));
   OAI21_X1 U2546 (.A(n340),
	.B1(n4021),
	.B2(n100),
	.ZN(n1362));
   NAND2_X1 U2547 (.A1(REGISTERS[255]),
	.A2(n4021),
	.ZN(n340));
   OAI21_X1 U2548 (.A(n406),
	.B1(FE_OFN80_n4035),
	.B2(n96),
	.ZN(n1424));
   NAND2_X1 U2549 (.A1(REGISTERS[317]),
	.A2(FE_OFN80_n4035),
	.ZN(n406));
   OAI21_X1 U2550 (.A(n407),
	.B1(FE_OFN80_n4035),
	.B2(n98),
	.ZN(n1425));
   NAND2_X1 U2551 (.A1(REGISTERS[318]),
	.A2(FE_OFN80_n4035),
	.ZN(n407));
   OAI21_X1 U2552 (.A(n439),
	.B1(FE_OFN59_n4034),
	.B2(n96),
	.ZN(n1456));
   NAND2_X1 U2553 (.A1(REGISTERS[349]),
	.A2(FE_OFN59_n4034),
	.ZN(n439));
   OAI21_X1 U2554 (.A(n440),
	.B1(FE_OFN59_n4034),
	.B2(n98),
	.ZN(n1457));
   NAND2_X1 U2555 (.A1(REGISTERS[350]),
	.A2(FE_OFN59_n4034),
	.ZN(n440));
   OAI21_X1 U2556 (.A(n472),
	.B1(FE_OFN70_n4033),
	.B2(n96),
	.ZN(n1488));
   NAND2_X1 U2557 (.A1(REGISTERS[381]),
	.A2(FE_OFN70_n4033),
	.ZN(n472));
   OAI21_X1 U2558 (.A(n473),
	.B1(FE_OFN70_n4033),
	.B2(n98),
	.ZN(n1489));
   NAND2_X1 U2559 (.A1(REGISTERS[382]),
	.A2(FE_OFN70_n4033),
	.ZN(n473));
   OAI21_X1 U2560 (.A(n505),
	.B1(FE_OFN87_n4032),
	.B2(n96),
	.ZN(n1520));
   NAND2_X1 U2561 (.A1(REGISTERS[413]),
	.A2(FE_OFN87_n4032),
	.ZN(n505));
   OAI21_X1 U2562 (.A(n506),
	.B1(FE_OFN87_n4032),
	.B2(n98),
	.ZN(n1521));
   NAND2_X1 U2563 (.A1(REGISTERS[414]),
	.A2(FE_OFN87_n4032),
	.ZN(n506));
   OAI21_X1 U2564 (.A(n538),
	.B1(FE_OFN63_n4031),
	.B2(n96),
	.ZN(n1552));
   NAND2_X1 U2565 (.A1(REGISTERS[445]),
	.A2(FE_OFN63_n4031),
	.ZN(n538));
   OAI21_X1 U2566 (.A(n539),
	.B1(FE_OFN63_n4031),
	.B2(n98),
	.ZN(n1553));
   NAND2_X1 U2567 (.A1(REGISTERS[446]),
	.A2(FE_OFN63_n4031),
	.ZN(n539));
   OAI21_X1 U2568 (.A(n571),
	.B1(FE_OFN81_n4030),
	.B2(n96),
	.ZN(n1584));
   NAND2_X1 U2569 (.A1(REGISTERS[477]),
	.A2(FE_OFN81_n4030),
	.ZN(n571));
   OAI21_X1 U2570 (.A(n572),
	.B1(FE_OFN81_n4030),
	.B2(n98),
	.ZN(n1585));
   NAND2_X1 U2571 (.A1(REGISTERS[478]),
	.A2(FE_OFN81_n4030),
	.ZN(n572));
   OAI21_X1 U2572 (.A(n604),
	.B1(FE_OFN67_n4029),
	.B2(n96),
	.ZN(n1616));
   NAND2_X1 U2573 (.A1(REGISTERS[509]),
	.A2(FE_OFN67_n4029),
	.ZN(n604));
   OAI21_X1 U2574 (.A(n605),
	.B1(FE_OFN67_n4029),
	.B2(n98),
	.ZN(n1617));
   NAND2_X1 U2575 (.A1(REGISTERS[510]),
	.A2(FE_OFN67_n4029),
	.ZN(n605));
   OAI21_X1 U2576 (.A(n637),
	.B1(n4019),
	.B2(n96),
	.ZN(n1648));
   NAND2_X1 U2577 (.A1(REGISTERS[541]),
	.A2(n4019),
	.ZN(n637));
   OAI21_X1 U2578 (.A(n638),
	.B1(FE_OFN61_n4019),
	.B2(n98),
	.ZN(n1649));
   NAND2_X1 U2579 (.A1(REGISTERS[542]),
	.A2(FE_OFN61_n4019),
	.ZN(n638));
   OAI21_X1 U2580 (.A(n671),
	.B1(FE_OFN65_n4018),
	.B2(n96),
	.ZN(n1680));
   NAND2_X1 U2581 (.A1(REGISTERS[573]),
	.A2(FE_OFN65_n4018),
	.ZN(n671));
   OAI21_X1 U2582 (.A(n672),
	.B1(FE_OFN65_n4018),
	.B2(n98),
	.ZN(n1681));
   NAND2_X1 U2583 (.A1(REGISTERS[574]),
	.A2(FE_OFN65_n4018),
	.ZN(n672));
   OAI21_X1 U2584 (.A(n704),
	.B1(n4017),
	.B2(n96),
	.ZN(n1712));
   NAND2_X1 U2585 (.A1(REGISTERS[605]),
	.A2(n4017),
	.ZN(n704));
   OAI21_X1 U2586 (.A(n705),
	.B1(FE_OFN66_n4017),
	.B2(n98),
	.ZN(n1713));
   NAND2_X1 U2587 (.A1(REGISTERS[606]),
	.A2(FE_OFN66_n4017),
	.ZN(n705));
   OAI21_X1 U2588 (.A(n737),
	.B1(FE_OFN62_n4016),
	.B2(n96),
	.ZN(n1744));
   NAND2_X1 U2589 (.A1(REGISTERS[637]),
	.A2(FE_OFN62_n4016),
	.ZN(n737));
   OAI21_X1 U2590 (.A(n738),
	.B1(FE_OFN62_n4016),
	.B2(n98),
	.ZN(n1745));
   NAND2_X1 U2591 (.A1(REGISTERS[638]),
	.A2(FE_OFN62_n4016),
	.ZN(n738));
   OAI21_X1 U2592 (.A(n770),
	.B1(n4015),
	.B2(n96),
	.ZN(n1776));
   NAND2_X1 U2593 (.A1(REGISTERS[669]),
	.A2(n4015),
	.ZN(n770));
   OAI21_X1 U2594 (.A(n771),
	.B1(FE_OFN74_n4015),
	.B2(n98),
	.ZN(n1777));
   NAND2_X1 U2595 (.A1(REGISTERS[670]),
	.A2(FE_OFN74_n4015),
	.ZN(n771));
   OAI21_X1 U2596 (.A(n803),
	.B1(n4014),
	.B2(n96),
	.ZN(n1808));
   NAND2_X1 U2597 (.A1(REGISTERS[701]),
	.A2(n4014),
	.ZN(n803));
   OAI21_X1 U2598 (.A(n804),
	.B1(FE_OFN78_n4014),
	.B2(n98),
	.ZN(n1809));
   NAND2_X1 U2599 (.A1(REGISTERS[702]),
	.A2(FE_OFN78_n4014),
	.ZN(n804));
   OAI21_X1 U2600 (.A(n836),
	.B1(n4013),
	.B2(n96),
	.ZN(n1840));
   NAND2_X1 U2601 (.A1(REGISTERS[733]),
	.A2(n4013),
	.ZN(n836));
   OAI21_X1 U2602 (.A(n837),
	.B1(FE_OFN76_n4013),
	.B2(n98),
	.ZN(n1841));
   NAND2_X1 U2603 (.A1(REGISTERS[734]),
	.A2(FE_OFN76_n4013),
	.ZN(n837));
   OAI21_X1 U2604 (.A(n869),
	.B1(n4012),
	.B2(n96),
	.ZN(n1872));
   NAND2_X1 U2605 (.A1(REGISTERS[765]),
	.A2(n4012),
	.ZN(n869));
   OAI21_X1 U2606 (.A(n870),
	.B1(FE_OFN64_n4012),
	.B2(n98),
	.ZN(n1873));
   NAND2_X1 U2607 (.A1(REGISTERS[766]),
	.A2(FE_OFN64_n4012),
	.ZN(n870));
   OAI21_X1 U2608 (.A(n1072),
	.B1(n4005),
	.B2(n38),
	.ZN(n2067));
   NAND2_X1 U2609 (.A1(REGISTERS[960]),
	.A2(n4005),
	.ZN(n1072));
   OAI21_X1 U2610 (.A(n1073),
	.B1(n4005),
	.B2(n40),
	.ZN(n2068));
   NAND2_X1 U2611 (.A1(REGISTERS[961]),
	.A2(n4005),
	.ZN(n1073));
   OAI21_X1 U2612 (.A(n1074),
	.B1(FE_OFN84_n4005),
	.B2(n42),
	.ZN(n2069));
   NAND2_X1 U2613 (.A1(REGISTERS[962]),
	.A2(FE_OFN84_n4005),
	.ZN(n1074));
   OAI21_X1 U2614 (.A(n1075),
	.B1(FE_OFN84_n4005),
	.B2(n44),
	.ZN(n2070));
   NAND2_X1 U2615 (.A1(REGISTERS[963]),
	.A2(FE_OFN84_n4005),
	.ZN(n1075));
   OAI21_X1 U2616 (.A(n1076),
	.B1(FE_OFN84_n4005),
	.B2(n46),
	.ZN(n2071));
   NAND2_X1 U2617 (.A1(REGISTERS[964]),
	.A2(FE_OFN84_n4005),
	.ZN(n1076));
   OAI21_X1 U2618 (.A(n1077),
	.B1(FE_OFN84_n4005),
	.B2(n48),
	.ZN(n2072));
   NAND2_X1 U2619 (.A1(REGISTERS[965]),
	.A2(FE_OFN84_n4005),
	.ZN(n1077));
   OAI21_X1 U2620 (.A(n1078),
	.B1(n4005),
	.B2(n50),
	.ZN(n2073));
   NAND2_X1 U2621 (.A1(REGISTERS[966]),
	.A2(n4005),
	.ZN(n1078));
   OAI21_X1 U2622 (.A(n1085),
	.B1(n4005),
	.B2(n64),
	.ZN(n2080));
   NAND2_X1 U2623 (.A1(REGISTERS[973]),
	.A2(n4005),
	.ZN(n1085));
   OAI21_X1 U2624 (.A(n1088),
	.B1(FE_OFN84_n4005),
	.B2(n70),
	.ZN(n2083));
   NAND2_X1 U2625 (.A1(REGISTERS[976]),
	.A2(FE_OFN84_n4005),
	.ZN(n1088));
   OAI21_X1 U2626 (.A(n1089),
	.B1(FE_OFN84_n4005),
	.B2(n72),
	.ZN(n2084));
   NAND2_X1 U2627 (.A1(REGISTERS[977]),
	.A2(FE_OFN84_n4005),
	.ZN(n1089));
   OAI21_X1 U2628 (.A(n1090),
	.B1(n4005),
	.B2(n74),
	.ZN(n2085));
   NAND2_X1 U2629 (.A1(REGISTERS[978]),
	.A2(n4005),
	.ZN(n1090));
   OAI21_X1 U2630 (.A(n1091),
	.B1(FE_OFN84_n4005),
	.B2(n76),
	.ZN(n2086));
   NAND2_X1 U2631 (.A1(REGISTERS[979]),
	.A2(FE_OFN84_n4005),
	.ZN(n1091));
   OAI21_X1 U2632 (.A(n1092),
	.B1(n4005),
	.B2(n78),
	.ZN(n2087));
   NAND2_X1 U2633 (.A1(REGISTERS[980]),
	.A2(n4005),
	.ZN(n1092));
   OAI21_X1 U2634 (.A(n1093),
	.B1(FE_OFN84_n4005),
	.B2(n80),
	.ZN(n2088));
   NAND2_X1 U2635 (.A1(REGISTERS[981]),
	.A2(FE_OFN84_n4005),
	.ZN(n1093));
   OAI21_X1 U2636 (.A(n1094),
	.B1(FE_OFN84_n4005),
	.B2(n82),
	.ZN(n2089));
   NAND2_X1 U2637 (.A1(REGISTERS[982]),
	.A2(FE_OFN84_n4005),
	.ZN(n1094));
   OAI21_X1 U2638 (.A(n1095),
	.B1(FE_OFN84_n4005),
	.B2(n84),
	.ZN(n2090));
   NAND2_X1 U2639 (.A1(REGISTERS[983]),
	.A2(FE_OFN84_n4005),
	.ZN(n1095));
   OAI21_X1 U2640 (.A(n1096),
	.B1(n4005),
	.B2(n86),
	.ZN(n2091));
   NAND2_X1 U2641 (.A1(REGISTERS[984]),
	.A2(n4005),
	.ZN(n1096));
   OAI21_X1 U2642 (.A(n1097),
	.B1(FE_OFN84_n4005),
	.B2(n88),
	.ZN(n2092));
   NAND2_X1 U2643 (.A1(REGISTERS[985]),
	.A2(FE_OFN84_n4005),
	.ZN(n1097));
   OAI21_X1 U2644 (.A(n1098),
	.B1(n4005),
	.B2(n90),
	.ZN(n2093));
   NAND2_X1 U2645 (.A1(REGISTERS[986]),
	.A2(n4005),
	.ZN(n1098));
   OAI21_X1 U2646 (.A(n1099),
	.B1(FE_OFN84_n4005),
	.B2(n92),
	.ZN(n2094));
   NAND2_X1 U2647 (.A1(REGISTERS[987]),
	.A2(FE_OFN84_n4005),
	.ZN(n1099));
   OAI21_X1 U2648 (.A(n1100),
	.B1(FE_OFN84_n4005),
	.B2(n94),
	.ZN(n2095));
   NAND2_X1 U2649 (.A1(REGISTERS[988]),
	.A2(FE_OFN84_n4005),
	.ZN(n1100));
   OAI21_X1 U2650 (.A(n1103),
	.B1(n4005),
	.B2(n100),
	.ZN(n2098));
   NAND2_X1 U2651 (.A1(REGISTERS[991]),
	.A2(n4005),
	.ZN(n1103));
   AND2_X1 U2652 (.A1(REGISTERS[992]),
	.A2(n4041),
	.ZN(n2099));
   AND2_X1 U2653 (.A1(REGISTERS[993]),
	.A2(n4041),
	.ZN(n2100));
   AND2_X1 U2654 (.A1(REGISTERS[994]),
	.A2(FE_OFN18_n4041),
	.ZN(n2101));
   AND2_X1 U2655 (.A1(REGISTERS[995]),
	.A2(FE_OFN18_n4041),
	.ZN(n2102));
   AND2_X1 U2656 (.A1(REGISTERS[996]),
	.A2(FE_OFN18_n4041),
	.ZN(n2103));
   AND2_X1 U2657 (.A1(REGISTERS[997]),
	.A2(FE_OFN18_n4041),
	.ZN(n2104));
   AND2_X1 U2658 (.A1(REGISTERS[998]),
	.A2(n4041),
	.ZN(n2105));
   AND2_X1 U2659 (.A1(REGISTERS[999]),
	.A2(FE_OFN18_n4041),
	.ZN(n2106));
   AND2_X1 U2660 (.A1(REGISTERS[1000]),
	.A2(n4041),
	.ZN(n2107));
   AND2_X1 U2661 (.A1(REGISTERS[1001]),
	.A2(FE_OFN18_n4041),
	.ZN(n2108));
   AND2_X1 U2662 (.A1(REGISTERS[1002]),
	.A2(n4041),
	.ZN(n2109));
   AND2_X1 U2663 (.A1(REGISTERS[1003]),
	.A2(FE_OFN18_n4041),
	.ZN(n2110));
   AND2_X1 U2664 (.A1(REGISTERS[1004]),
	.A2(n4041),
	.ZN(n2111));
   AND2_X1 U2665 (.A1(REGISTERS[1005]),
	.A2(n4041),
	.ZN(n2112));
   AND2_X1 U2666 (.A1(REGISTERS[1006]),
	.A2(FE_OFN18_n4041),
	.ZN(n2113));
   AND2_X1 U2667 (.A1(REGISTERS[1007]),
	.A2(FE_OFN18_n4041),
	.ZN(n2114));
   AND2_X1 U2668 (.A1(REGISTERS[1008]),
	.A2(FE_OFN18_n4041),
	.ZN(n2115));
   AND2_X1 U2669 (.A1(REGISTERS[1009]),
	.A2(FE_OFN18_n4041),
	.ZN(n2116));
   AND2_X1 U2670 (.A1(REGISTERS[1010]),
	.A2(n4041),
	.ZN(n2117));
   AND2_X1 U2671 (.A1(REGISTERS[1011]),
	.A2(FE_OFN18_n4041),
	.ZN(n2118));
   AND2_X1 U2672 (.A1(REGISTERS[1012]),
	.A2(n4041),
	.ZN(n2119));
   AND2_X1 U2673 (.A1(REGISTERS[1013]),
	.A2(FE_OFN18_n4041),
	.ZN(n2120));
   AND2_X1 U2674 (.A1(REGISTERS[1014]),
	.A2(FE_OFN18_n4041),
	.ZN(n2121));
   AND2_X1 U2675 (.A1(REGISTERS[1015]),
	.A2(FE_OFN18_n4041),
	.ZN(n2122));
   AND2_X1 U2676 (.A1(REGISTERS[1016]),
	.A2(n4041),
	.ZN(n2123));
   AND2_X1 U2677 (.A1(REGISTERS[1017]),
	.A2(FE_OFN18_n4041),
	.ZN(n2124));
   AND2_X1 U2678 (.A1(REGISTERS[1018]),
	.A2(n4041),
	.ZN(n2125));
   AND2_X1 U2679 (.A1(REGISTERS[1019]),
	.A2(FE_OFN18_n4041),
	.ZN(n2126));
   AND2_X1 U2680 (.A1(REGISTERS[1020]),
	.A2(FE_OFN18_n4041),
	.ZN(n2127));
   AND2_X1 U2681 (.A1(REGISTERS[1021]),
	.A2(n4041),
	.ZN(n2128));
   AND2_X1 U2682 (.A1(REGISTERS[1022]),
	.A2(FE_OFN18_n4041),
	.ZN(n2129));
   AND2_X1 U2683 (.A1(REGISTERS[1023]),
	.A2(n4041),
	.ZN(n2130));
   NAND2_X2 U2684 (.A1(ADD_RD1[4]),
	.A2(n2785),
	.ZN(n2780));
   NOR2_X1 U2685 (.A1(n2784),
	.A2(ADD_RD1[1]),
	.ZN(n1));
   AND2_X2 U2686 (.A1(n1),
	.A2(ADD_RD1[0]),
	.ZN(n2762));
   NOR2_X1 U2687 (.A1(n2784),
	.A2(n2783),
	.ZN(n2));
   AND2_X2 U2688 (.A1(ADD_RD1[0]),
	.A2(n2),
	.ZN(n2761));
   AOI22_X1 U2689 (.A1(REGISTERS[320]),
	.A2(FE_OFN13_n2762),
	.B1(REGISTERS[256]),
	.B2(FE_OFN135_n2761),
	.ZN(n8));
   NOR2_X1 U2690 (.A1(ADD_RD1[1]),
	.A2(ADD_RD1[2]),
	.ZN(n3));
   AND2_X2 U2691 (.A1(n3),
	.A2(ADD_RD1[0]),
	.ZN(n2764));
   NOR2_X1 U2692 (.A1(n2783),
	.A2(ADD_RD1[2]),
	.ZN(n4));
   AND2_X2 U2693 (.A1(n4),
	.A2(ADD_RD1[0]),
	.ZN(n2763));
   AOI22_X1 U2694 (.A1(REGISTERS[448]),
	.A2(FE_OFN54_n2764),
	.B1(REGISTERS[384]),
	.B2(FE_OFN110_n2763),
	.ZN(n7));
   AND2_X1 U2695 (.A1(n1),
	.A2(n2782),
	.ZN(n2766));
   AND2_X2 U2696 (.A1(n2),
	.A2(n2782),
	.ZN(n2765));
   AOI22_X1 U2697 (.A1(REGISTERS[352]),
	.A2(FE_OFN9_n2766),
	.B1(REGISTERS[288]),
	.B2(n2765),
	.ZN(n6));
   AND2_X2 U2698 (.A1(n3),
	.A2(n2782),
	.ZN(n2768));
   AND2_X2 U2699 (.A1(n4),
	.A2(n2782),
	.ZN(n2767));
   AOI22_X1 U2700 (.A1(REGISTERS[480]),
	.A2(n2768),
	.B1(REGISTERS[416]),
	.B2(n2767),
	.ZN(n5));
   AND4_X1 U2701 (.A1(n8),
	.A2(n7),
	.A3(n6),
	.A4(n5),
	.ZN(n25));
   NAND2_X2 U2702 (.A1(ADD_RD1[4]),
	.A2(ADD_RD1[3]),
	.ZN(n2778));
   AOI22_X1 U2703 (.A1(REGISTERS[64]),
	.A2(FE_OFN13_n2762),
	.B1(REGISTERS[0]),
	.B2(FE_OFN135_n2761),
	.ZN(n12));
   AOI22_X1 U2704 (.A1(REGISTERS[192]),
	.A2(FE_OFN54_n2764),
	.B1(REGISTERS[128]),
	.B2(FE_OFN110_n2763),
	.ZN(n11));
   AOI22_X1 U2705 (.A1(REGISTERS[96]),
	.A2(FE_OFN9_n2766),
	.B1(REGISTERS[32]),
	.B2(n2765),
	.ZN(n10));
   AOI22_X1 U2706 (.A1(REGISTERS[224]),
	.A2(n2768),
	.B1(REGISTERS[160]),
	.B2(n2767),
	.ZN(n9));
   AND4_X1 U2707 (.A1(n12),
	.A2(n11),
	.A3(n10),
	.A4(n9),
	.ZN(n24));
   AOI22_X1 U2708 (.A1(REGISTERS[832]),
	.A2(n2762),
	.B1(REGISTERS[768]),
	.B2(n2761),
	.ZN(n16));
   AOI22_X1 U2709 (.A1(REGISTERS[960]),
	.A2(FE_OFN54_n2764),
	.B1(REGISTERS[896]),
	.B2(FE_OFN110_n2763),
	.ZN(n15));
   AOI22_X1 U2710 (.A1(REGISTERS[864]),
	.A2(FE_OFN9_n2766),
	.B1(REGISTERS[800]),
	.B2(n2765),
	.ZN(n14));
   AOI22_X1 U2711 (.A1(REGISTERS[992]),
	.A2(n2768),
	.B1(REGISTERS[928]),
	.B2(n2767),
	.ZN(n13));
   NAND4_X1 U2712 (.A1(n16),
	.A2(n15),
	.A3(n14),
	.A4(n13),
	.ZN(n22));
   NOR2_X1 U2713 (.A1(ADD_RD1[3]),
	.A2(ADD_RD1[4]),
	.ZN(n2776));
   AOI22_X1 U2714 (.A1(REGISTERS[576]),
	.A2(n2762),
	.B1(REGISTERS[512]),
	.B2(n2761),
	.ZN(n20));
   AOI22_X1 U2715 (.A1(REGISTERS[704]),
	.A2(FE_OFN54_n2764),
	.B1(REGISTERS[640]),
	.B2(FE_OFN110_n2763),
	.ZN(n19));
   AOI22_X1 U2716 (.A1(REGISTERS[608]),
	.A2(FE_OFN9_n2766),
	.B1(REGISTERS[544]),
	.B2(n2765),
	.ZN(n18));
   AOI22_X1 U2717 (.A1(REGISTERS[736]),
	.A2(n2768),
	.B1(REGISTERS[672]),
	.B2(n2767),
	.ZN(n17));
   NAND4_X1 U2718 (.A1(n20),
	.A2(n19),
	.A3(n18),
	.A4(n17),
	.ZN(n21));
   NOR2_X1 U2719 (.A1(n2785),
	.A2(ADD_RD1[4]),
	.ZN(n2774));
   AOI22_X1 U2720 (.A1(n22),
	.A2(FE_OFN32_n2776),
	.B1(n21),
	.B2(FE_OFN30_n2774),
	.ZN(n23));
   OAI221_X1 U2721 (.A(n23),
	.B1(n2780),
	.B2(n25),
	.C1(n2778),
	.C2(n24),
	.ZN(N62));
   AOI22_X1 U2722 (.A1(REGISTERS[321]),
	.A2(FE_OFN13_n2762),
	.B1(REGISTERS[257]),
	.B2(FE_OFN135_n2761),
	.ZN(n29));
   AOI22_X1 U2723 (.A1(REGISTERS[449]),
	.A2(n2764),
	.B1(REGISTERS[385]),
	.B2(n2763),
	.ZN(n28));
   AOI22_X1 U2724 (.A1(REGISTERS[353]),
	.A2(FE_OFN8_n2766),
	.B1(REGISTERS[289]),
	.B2(FE_OFN51_n2765),
	.ZN(n27));
   AOI22_X1 U2725 (.A1(REGISTERS[481]),
	.A2(FE_OFN113_n2768),
	.B1(REGISTERS[417]),
	.B2(FE_OFN11_n2767),
	.ZN(n26));
   AND4_X1 U2726 (.A1(n29),
	.A2(n28),
	.A3(n27),
	.A4(n26),
	.ZN(n2139));
   AOI22_X1 U2727 (.A1(REGISTERS[65]),
	.A2(FE_OFN13_n2762),
	.B1(REGISTERS[1]),
	.B2(FE_OFN135_n2761),
	.ZN(n33));
   AOI22_X1 U2728 (.A1(REGISTERS[193]),
	.A2(n2764),
	.B1(REGISTERS[129]),
	.B2(n2763),
	.ZN(n32));
   AOI22_X1 U2729 (.A1(REGISTERS[97]),
	.A2(FE_OFN8_n2766),
	.B1(REGISTERS[33]),
	.B2(FE_OFN51_n2765),
	.ZN(n31));
   AOI22_X1 U2730 (.A1(REGISTERS[225]),
	.A2(FE_OFN113_n2768),
	.B1(REGISTERS[161]),
	.B2(FE_OFN11_n2767),
	.ZN(n30));
   AND4_X1 U2731 (.A1(n33),
	.A2(n32),
	.A3(n31),
	.A4(n30),
	.ZN(n2138));
   AOI22_X1 U2732 (.A1(REGISTERS[833]),
	.A2(FE_OFN13_n2762),
	.B1(REGISTERS[769]),
	.B2(FE_OFN135_n2761),
	.ZN(n37));
   AOI22_X1 U2733 (.A1(REGISTERS[961]),
	.A2(FE_OFN54_n2764),
	.B1(REGISTERS[897]),
	.B2(FE_OFN110_n2763),
	.ZN(n36));
   AOI22_X1 U2734 (.A1(REGISTERS[865]),
	.A2(FE_OFN8_n2766),
	.B1(REGISTERS[801]),
	.B2(n2765),
	.ZN(n35));
   AOI22_X1 U2735 (.A1(REGISTERS[993]),
	.A2(FE_OFN113_n2768),
	.B1(REGISTERS[929]),
	.B2(FE_OFN11_n2767),
	.ZN(n34));
   NAND4_X1 U2736 (.A1(n37),
	.A2(n36),
	.A3(n35),
	.A4(n34),
	.ZN(n2136));
   AOI22_X1 U2737 (.A1(REGISTERS[577]),
	.A2(FE_OFN13_n2762),
	.B1(REGISTERS[513]),
	.B2(FE_OFN135_n2761),
	.ZN(n2134));
   AOI22_X1 U2738 (.A1(REGISTERS[705]),
	.A2(FE_OFN54_n2764),
	.B1(REGISTERS[641]),
	.B2(FE_OFN110_n2763),
	.ZN(n2133));
   AOI22_X1 U2739 (.A1(REGISTERS[609]),
	.A2(FE_OFN8_n2766),
	.B1(REGISTERS[545]),
	.B2(n2765),
	.ZN(n2132));
   AOI22_X1 U2740 (.A1(REGISTERS[737]),
	.A2(FE_OFN113_n2768),
	.B1(REGISTERS[673]),
	.B2(FE_OFN11_n2767),
	.ZN(n2131));
   NAND4_X1 U2741 (.A1(n2134),
	.A2(n2133),
	.A3(n2132),
	.A4(n2131),
	.ZN(n2135));
   AOI22_X1 U2742 (.A1(n2136),
	.A2(FE_OFN32_n2776),
	.B1(n2135),
	.B2(FE_OFN30_n2774),
	.ZN(n2137));
   OAI221_X1 U2743 (.A(n2137),
	.B1(n2780),
	.B2(n2139),
	.C1(n2778),
	.C2(n2138),
	.ZN(N61));
   AOI22_X1 U2744 (.A1(REGISTERS[322]),
	.A2(FE_OFN13_n2762),
	.B1(REGISTERS[258]),
	.B2(FE_OFN135_n2761),
	.ZN(n2143));
   AOI22_X1 U2745 (.A1(REGISTERS[450]),
	.A2(FE_OFN55_n2764),
	.B1(REGISTERS[386]),
	.B2(FE_OFN111_n2763),
	.ZN(n2142));
   AOI22_X1 U2746 (.A1(REGISTERS[354]),
	.A2(FE_OFN9_n2766),
	.B1(REGISTERS[290]),
	.B2(n2765),
	.ZN(n2141));
   AOI22_X1 U2747 (.A1(REGISTERS[482]),
	.A2(FE_OFN113_n2768),
	.B1(REGISTERS[418]),
	.B2(FE_OFN11_n2767),
	.ZN(n2140));
   AND4_X1 U2748 (.A1(n2143),
	.A2(n2142),
	.A3(n2141),
	.A4(n2140),
	.ZN(n2160));
   AOI22_X1 U2749 (.A1(REGISTERS[66]),
	.A2(FE_OFN13_n2762),
	.B1(REGISTERS[2]),
	.B2(FE_OFN135_n2761),
	.ZN(n2147));
   AOI22_X1 U2750 (.A1(REGISTERS[194]),
	.A2(FE_OFN55_n2764),
	.B1(REGISTERS[130]),
	.B2(FE_OFN111_n2763),
	.ZN(n2146));
   AOI22_X1 U2751 (.A1(REGISTERS[98]),
	.A2(FE_OFN9_n2766),
	.B1(REGISTERS[34]),
	.B2(n2765),
	.ZN(n2145));
   AOI22_X1 U2752 (.A1(REGISTERS[226]),
	.A2(FE_OFN113_n2768),
	.B1(REGISTERS[162]),
	.B2(FE_OFN11_n2767),
	.ZN(n2144));
   AND4_X1 U2753 (.A1(n2147),
	.A2(n2146),
	.A3(n2145),
	.A4(n2144),
	.ZN(n2159));
   AOI22_X1 U2754 (.A1(REGISTERS[834]),
	.A2(FE_OFN14_n2762),
	.B1(REGISTERS[770]),
	.B2(FE_OFN136_n2761),
	.ZN(n2151));
   AOI22_X1 U2755 (.A1(REGISTERS[962]),
	.A2(FE_OFN56_n2764),
	.B1(REGISTERS[898]),
	.B2(FE_OFN112_n2763),
	.ZN(n2150));
   AOI22_X1 U2756 (.A1(REGISTERS[866]),
	.A2(FE_OFN10_n2766),
	.B1(REGISTERS[802]),
	.B2(FE_OFN53_n2765),
	.ZN(n2149));
   AOI22_X1 U2757 (.A1(REGISTERS[994]),
	.A2(FE_OFN114_n2768),
	.B1(REGISTERS[930]),
	.B2(FE_OFN12_n2767),
	.ZN(n2148));
   NAND4_X1 U2758 (.A1(n2151),
	.A2(n2150),
	.A3(n2149),
	.A4(n2148),
	.ZN(n2157));
   AOI22_X1 U2759 (.A1(REGISTERS[578]),
	.A2(FE_OFN14_n2762),
	.B1(REGISTERS[514]),
	.B2(FE_OFN136_n2761),
	.ZN(n2155));
   AOI22_X1 U2760 (.A1(REGISTERS[706]),
	.A2(FE_OFN56_n2764),
	.B1(REGISTERS[642]),
	.B2(FE_OFN112_n2763),
	.ZN(n2154));
   AOI22_X1 U2761 (.A1(REGISTERS[610]),
	.A2(FE_OFN10_n2766),
	.B1(REGISTERS[546]),
	.B2(FE_OFN53_n2765),
	.ZN(n2153));
   AOI22_X1 U2762 (.A1(REGISTERS[738]),
	.A2(FE_OFN114_n2768),
	.B1(REGISTERS[674]),
	.B2(FE_OFN12_n2767),
	.ZN(n2152));
   NAND4_X1 U2763 (.A1(n2155),
	.A2(n2154),
	.A3(n2153),
	.A4(n2152),
	.ZN(n2156));
   AOI22_X1 U2764 (.A1(n2157),
	.A2(FE_OFN32_n2776),
	.B1(n2156),
	.B2(FE_OFN30_n2774),
	.ZN(n2158));
   OAI221_X1 U2765 (.A(n2158),
	.B1(n2780),
	.B2(n2160),
	.C1(n2778),
	.C2(n2159),
	.ZN(N60));
   AOI22_X1 U2766 (.A1(REGISTERS[323]),
	.A2(FE_OFN14_n2762),
	.B1(REGISTERS[259]),
	.B2(FE_OFN136_n2761),
	.ZN(n2164));
   AOI22_X1 U2767 (.A1(REGISTERS[451]),
	.A2(FE_OFN55_n2764),
	.B1(REGISTERS[387]),
	.B2(FE_OFN111_n2763),
	.ZN(n2163));
   AOI22_X1 U2768 (.A1(REGISTERS[355]),
	.A2(FE_OFN9_n2766),
	.B1(REGISTERS[291]),
	.B2(FE_OFN52_n2765),
	.ZN(n2162));
   AOI22_X1 U2769 (.A1(REGISTERS[483]),
	.A2(FE_OFN114_n2768),
	.B1(REGISTERS[419]),
	.B2(FE_OFN12_n2767),
	.ZN(n2161));
   AND4_X1 U2770 (.A1(n2164),
	.A2(n2163),
	.A3(n2162),
	.A4(n2161),
	.ZN(n2181));
   AOI22_X1 U2771 (.A1(REGISTERS[67]),
	.A2(FE_OFN14_n2762),
	.B1(REGISTERS[3]),
	.B2(FE_OFN136_n2761),
	.ZN(n2168));
   AOI22_X1 U2772 (.A1(REGISTERS[195]),
	.A2(FE_OFN55_n2764),
	.B1(REGISTERS[131]),
	.B2(FE_OFN111_n2763),
	.ZN(n2167));
   AOI22_X1 U2773 (.A1(REGISTERS[99]),
	.A2(FE_OFN9_n2766),
	.B1(REGISTERS[35]),
	.B2(FE_OFN52_n2765),
	.ZN(n2166));
   AOI22_X1 U2774 (.A1(REGISTERS[227]),
	.A2(FE_OFN114_n2768),
	.B1(REGISTERS[163]),
	.B2(FE_OFN12_n2767),
	.ZN(n2165));
   AND4_X1 U2775 (.A1(n2168),
	.A2(n2167),
	.A3(n2166),
	.A4(n2165),
	.ZN(n2180));
   AOI22_X1 U2776 (.A1(REGISTERS[835]),
	.A2(FE_OFN14_n2762),
	.B1(REGISTERS[771]),
	.B2(n2761),
	.ZN(n2172));
   AOI22_X1 U2777 (.A1(REGISTERS[963]),
	.A2(FE_OFN56_n2764),
	.B1(REGISTERS[899]),
	.B2(FE_OFN112_n2763),
	.ZN(n2171));
   AOI22_X1 U2778 (.A1(REGISTERS[867]),
	.A2(FE_OFN10_n2766),
	.B1(REGISTERS[803]),
	.B2(FE_OFN53_n2765),
	.ZN(n2170));
   AOI22_X1 U2779 (.A1(REGISTERS[995]),
	.A2(FE_OFN114_n2768),
	.B1(REGISTERS[931]),
	.B2(FE_OFN12_n2767),
	.ZN(n2169));
   NAND4_X1 U2780 (.A1(n2172),
	.A2(n2171),
	.A3(n2170),
	.A4(n2169),
	.ZN(n2178));
   AOI22_X1 U2781 (.A1(REGISTERS[579]),
	.A2(FE_OFN14_n2762),
	.B1(REGISTERS[515]),
	.B2(FE_OFN136_n2761),
	.ZN(n2176));
   AOI22_X1 U2782 (.A1(REGISTERS[707]),
	.A2(FE_OFN56_n2764),
	.B1(REGISTERS[643]),
	.B2(FE_OFN112_n2763),
	.ZN(n2175));
   AOI22_X1 U2783 (.A1(REGISTERS[611]),
	.A2(FE_OFN10_n2766),
	.B1(REGISTERS[547]),
	.B2(FE_OFN53_n2765),
	.ZN(n2174));
   AOI22_X1 U2784 (.A1(REGISTERS[739]),
	.A2(FE_OFN114_n2768),
	.B1(REGISTERS[675]),
	.B2(FE_OFN12_n2767),
	.ZN(n2173));
   NAND4_X1 U2785 (.A1(n2176),
	.A2(n2175),
	.A3(n2174),
	.A4(n2173),
	.ZN(n2177));
   AOI22_X1 U2786 (.A1(n2178),
	.A2(FE_OFN32_n2776),
	.B1(n2177),
	.B2(FE_OFN30_n2774),
	.ZN(n2179));
   OAI221_X1 U2787 (.A(n2179),
	.B1(n2780),
	.B2(n2181),
	.C1(n2778),
	.C2(n2180),
	.ZN(N59));
   AOI22_X1 U2788 (.A1(REGISTERS[324]),
	.A2(n2762),
	.B1(REGISTERS[260]),
	.B2(n2761),
	.ZN(n2185));
   AOI22_X1 U2789 (.A1(REGISTERS[452]),
	.A2(n2764),
	.B1(REGISTERS[388]),
	.B2(n2763),
	.ZN(n2184));
   AOI22_X1 U2790 (.A1(REGISTERS[356]),
	.A2(n2766),
	.B1(REGISTERS[292]),
	.B2(n2765),
	.ZN(n2183));
   AOI22_X1 U2791 (.A1(REGISTERS[484]),
	.A2(n2768),
	.B1(REGISTERS[420]),
	.B2(n2767),
	.ZN(n2182));
   AND4_X1 U2792 (.A1(n2185),
	.A2(n2184),
	.A3(n2183),
	.A4(n2182),
	.ZN(n2202));
   AOI22_X1 U2793 (.A1(REGISTERS[68]),
	.A2(n2762),
	.B1(REGISTERS[4]),
	.B2(n2761),
	.ZN(n2189));
   AOI22_X1 U2794 (.A1(REGISTERS[196]),
	.A2(n2764),
	.B1(REGISTERS[132]),
	.B2(n2763),
	.ZN(n2188));
   AOI22_X1 U2795 (.A1(REGISTERS[100]),
	.A2(FE_OFN8_n2766),
	.B1(REGISTERS[36]),
	.B2(n2765),
	.ZN(n2187));
   AOI22_X1 U2796 (.A1(REGISTERS[228]),
	.A2(n2768),
	.B1(REGISTERS[164]),
	.B2(n2767),
	.ZN(n2186));
   AND4_X1 U2797 (.A1(n2189),
	.A2(n2188),
	.A3(n2187),
	.A4(n2186),
	.ZN(n2201));
   AOI22_X1 U2798 (.A1(REGISTERS[836]),
	.A2(n2762),
	.B1(REGISTERS[772]),
	.B2(n2761),
	.ZN(n2193));
   AOI22_X1 U2799 (.A1(REGISTERS[964]),
	.A2(FE_OFN54_n2764),
	.B1(REGISTERS[900]),
	.B2(n2763),
	.ZN(n2192));
   AOI22_X1 U2800 (.A1(REGISTERS[868]),
	.A2(n2766),
	.B1(REGISTERS[804]),
	.B2(n2765),
	.ZN(n2191));
   AOI22_X1 U2801 (.A1(REGISTERS[996]),
	.A2(n2768),
	.B1(REGISTERS[932]),
	.B2(n2767),
	.ZN(n2190));
   NAND4_X1 U2802 (.A1(n2193),
	.A2(n2192),
	.A3(n2191),
	.A4(n2190),
	.ZN(n2199));
   AOI22_X1 U2803 (.A1(REGISTERS[580]),
	.A2(n2762),
	.B1(REGISTERS[516]),
	.B2(n2761),
	.ZN(n2197));
   AOI22_X1 U2804 (.A1(REGISTERS[708]),
	.A2(FE_OFN54_n2764),
	.B1(REGISTERS[644]),
	.B2(n2763),
	.ZN(n2196));
   AOI22_X1 U2805 (.A1(REGISTERS[612]),
	.A2(n2766),
	.B1(REGISTERS[548]),
	.B2(n2765),
	.ZN(n2195));
   AOI22_X1 U2806 (.A1(REGISTERS[740]),
	.A2(n2768),
	.B1(REGISTERS[676]),
	.B2(n2767),
	.ZN(n2194));
   NAND4_X1 U2807 (.A1(n2197),
	.A2(n2196),
	.A3(n2195),
	.A4(n2194),
	.ZN(n2198));
   AOI22_X1 U2808 (.A1(n2199),
	.A2(FE_OFN32_n2776),
	.B1(n2198),
	.B2(FE_OFN30_n2774),
	.ZN(n2200));
   OAI221_X1 U2809 (.A(n2200),
	.B1(n2780),
	.B2(n2202),
	.C1(n2778),
	.C2(n2201),
	.ZN(N58));
   AOI22_X1 U2810 (.A1(REGISTERS[325]),
	.A2(FE_OFN14_n2762),
	.B1(REGISTERS[261]),
	.B2(FE_OFN136_n2761),
	.ZN(n2206));
   AOI22_X1 U2811 (.A1(REGISTERS[453]),
	.A2(FE_OFN55_n2764),
	.B1(REGISTERS[389]),
	.B2(FE_OFN111_n2763),
	.ZN(n2205));
   AOI22_X1 U2812 (.A1(REGISTERS[357]),
	.A2(FE_OFN9_n2766),
	.B1(REGISTERS[293]),
	.B2(FE_OFN53_n2765),
	.ZN(n2204));
   AOI22_X1 U2813 (.A1(REGISTERS[485]),
	.A2(FE_OFN114_n2768),
	.B1(REGISTERS[421]),
	.B2(FE_OFN12_n2767),
	.ZN(n2203));
   AND4_X1 U2814 (.A1(n2206),
	.A2(n2205),
	.A3(n2204),
	.A4(n2203),
	.ZN(n2223));
   AOI22_X1 U2815 (.A1(REGISTERS[69]),
	.A2(FE_OFN14_n2762),
	.B1(REGISTERS[5]),
	.B2(FE_OFN136_n2761),
	.ZN(n2210));
   AOI22_X1 U2816 (.A1(REGISTERS[197]),
	.A2(FE_OFN55_n2764),
	.B1(REGISTERS[133]),
	.B2(FE_OFN111_n2763),
	.ZN(n2209));
   AOI22_X1 U2817 (.A1(REGISTERS[101]),
	.A2(FE_OFN9_n2766),
	.B1(REGISTERS[37]),
	.B2(FE_OFN53_n2765),
	.ZN(n2208));
   AOI22_X1 U2818 (.A1(REGISTERS[229]),
	.A2(FE_OFN114_n2768),
	.B1(REGISTERS[165]),
	.B2(FE_OFN12_n2767),
	.ZN(n2207));
   AND4_X1 U2819 (.A1(n2210),
	.A2(n2209),
	.A3(n2208),
	.A4(n2207),
	.ZN(n2222));
   AOI22_X1 U2820 (.A1(REGISTERS[837]),
	.A2(n2762),
	.B1(REGISTERS[773]),
	.B2(n2761),
	.ZN(n2214));
   AOI22_X1 U2821 (.A1(REGISTERS[965]),
	.A2(FE_OFN56_n2764),
	.B1(REGISTERS[901]),
	.B2(FE_OFN112_n2763),
	.ZN(n2213));
   AOI22_X1 U2822 (.A1(REGISTERS[869]),
	.A2(FE_OFN9_n2766),
	.B1(REGISTERS[805]),
	.B2(FE_OFN53_n2765),
	.ZN(n2212));
   AOI22_X1 U2823 (.A1(REGISTERS[997]),
	.A2(FE_OFN114_n2768),
	.B1(REGISTERS[933]),
	.B2(FE_OFN12_n2767),
	.ZN(n2211));
   NAND4_X1 U2824 (.A1(n2214),
	.A2(n2213),
	.A3(n2212),
	.A4(n2211),
	.ZN(n2220));
   AOI22_X1 U2825 (.A1(REGISTERS[581]),
	.A2(FE_OFN14_n2762),
	.B1(REGISTERS[517]),
	.B2(n2761),
	.ZN(n2218));
   AOI22_X1 U2826 (.A1(REGISTERS[709]),
	.A2(FE_OFN56_n2764),
	.B1(REGISTERS[645]),
	.B2(FE_OFN112_n2763),
	.ZN(n2217));
   AOI22_X1 U2827 (.A1(REGISTERS[613]),
	.A2(FE_OFN9_n2766),
	.B1(REGISTERS[549]),
	.B2(FE_OFN53_n2765),
	.ZN(n2216));
   AOI22_X1 U2828 (.A1(REGISTERS[741]),
	.A2(FE_OFN114_n2768),
	.B1(REGISTERS[677]),
	.B2(FE_OFN12_n2767),
	.ZN(n2215));
   NAND4_X1 U2829 (.A1(n2218),
	.A2(n2217),
	.A3(n2216),
	.A4(n2215),
	.ZN(n2219));
   AOI22_X1 U2830 (.A1(n2220),
	.A2(FE_OFN32_n2776),
	.B1(n2219),
	.B2(FE_OFN30_n2774),
	.ZN(n2221));
   OAI221_X1 U2831 (.A(n2221),
	.B1(n2780),
	.B2(n2223),
	.C1(n2778),
	.C2(n2222),
	.ZN(N57));
   AOI22_X1 U2832 (.A1(REGISTERS[326]),
	.A2(FE_OFN13_n2762),
	.B1(REGISTERS[262]),
	.B2(FE_OFN135_n2761),
	.ZN(n2227));
   AOI22_X1 U2833 (.A1(REGISTERS[454]),
	.A2(n2764),
	.B1(REGISTERS[390]),
	.B2(n2763),
	.ZN(n2226));
   AOI22_X1 U2834 (.A1(REGISTERS[358]),
	.A2(FE_OFN8_n2766),
	.B1(REGISTERS[294]),
	.B2(FE_OFN51_n2765),
	.ZN(n2225));
   AOI22_X1 U2835 (.A1(REGISTERS[486]),
	.A2(FE_OFN113_n2768),
	.B1(REGISTERS[422]),
	.B2(n2767),
	.ZN(n2224));
   AND4_X1 U2836 (.A1(n2227),
	.A2(n2226),
	.A3(n2225),
	.A4(n2224),
	.ZN(n2244));
   AOI22_X1 U2837 (.A1(REGISTERS[70]),
	.A2(FE_OFN13_n2762),
	.B1(REGISTERS[6]),
	.B2(FE_OFN135_n2761),
	.ZN(n2231));
   AOI22_X1 U2838 (.A1(REGISTERS[198]),
	.A2(n2764),
	.B1(REGISTERS[134]),
	.B2(n2763),
	.ZN(n2230));
   AOI22_X1 U2839 (.A1(REGISTERS[102]),
	.A2(FE_OFN8_n2766),
	.B1(REGISTERS[38]),
	.B2(FE_OFN51_n2765),
	.ZN(n2229));
   AOI22_X1 U2840 (.A1(REGISTERS[230]),
	.A2(FE_OFN113_n2768),
	.B1(REGISTERS[166]),
	.B2(n2767),
	.ZN(n2228));
   AND4_X1 U2841 (.A1(n2231),
	.A2(n2230),
	.A3(n2229),
	.A4(n2228),
	.ZN(n2243));
   AOI22_X1 U2842 (.A1(REGISTERS[838]),
	.A2(FE_OFN13_n2762),
	.B1(REGISTERS[774]),
	.B2(FE_OFN135_n2761),
	.ZN(n2235));
   AOI22_X1 U2843 (.A1(REGISTERS[966]),
	.A2(FE_OFN54_n2764),
	.B1(REGISTERS[902]),
	.B2(FE_OFN110_n2763),
	.ZN(n2234));
   AOI22_X1 U2844 (.A1(REGISTERS[870]),
	.A2(FE_OFN8_n2766),
	.B1(REGISTERS[806]),
	.B2(n2765),
	.ZN(n2233));
   AOI22_X1 U2845 (.A1(REGISTERS[998]),
	.A2(FE_OFN113_n2768),
	.B1(REGISTERS[934]),
	.B2(FE_OFN11_n2767),
	.ZN(n2232));
   NAND4_X1 U2846 (.A1(n2235),
	.A2(n2234),
	.A3(n2233),
	.A4(n2232),
	.ZN(n2241));
   AOI22_X1 U2847 (.A1(REGISTERS[582]),
	.A2(FE_OFN13_n2762),
	.B1(REGISTERS[518]),
	.B2(FE_OFN135_n2761),
	.ZN(n2239));
   AOI22_X1 U2848 (.A1(REGISTERS[710]),
	.A2(FE_OFN54_n2764),
	.B1(REGISTERS[646]),
	.B2(FE_OFN110_n2763),
	.ZN(n2238));
   AOI22_X1 U2849 (.A1(REGISTERS[614]),
	.A2(FE_OFN9_n2766),
	.B1(REGISTERS[550]),
	.B2(n2765),
	.ZN(n2237));
   AOI22_X1 U2850 (.A1(REGISTERS[742]),
	.A2(FE_OFN113_n2768),
	.B1(REGISTERS[678]),
	.B2(FE_OFN11_n2767),
	.ZN(n2236));
   NAND4_X1 U2851 (.A1(n2239),
	.A2(n2238),
	.A3(n2237),
	.A4(n2236),
	.ZN(n2240));
   AOI22_X1 U2852 (.A1(n2241),
	.A2(FE_OFN32_n2776),
	.B1(n2240),
	.B2(FE_OFN30_n2774),
	.ZN(n2242));
   OAI221_X1 U2853 (.A(n2242),
	.B1(n2780),
	.B2(n2244),
	.C1(n2778),
	.C2(n2243),
	.ZN(N56));
   AOI22_X1 U2854 (.A1(REGISTERS[327]),
	.A2(FE_OFN14_n2762),
	.B1(REGISTERS[263]),
	.B2(FE_OFN136_n2761),
	.ZN(n2248));
   AOI22_X1 U2855 (.A1(REGISTERS[455]),
	.A2(FE_OFN55_n2764),
	.B1(REGISTERS[391]),
	.B2(FE_OFN111_n2763),
	.ZN(n2247));
   AOI22_X1 U2856 (.A1(REGISTERS[359]),
	.A2(FE_OFN9_n2766),
	.B1(REGISTERS[295]),
	.B2(FE_OFN52_n2765),
	.ZN(n2246));
   AOI22_X1 U2857 (.A1(REGISTERS[487]),
	.A2(FE_OFN114_n2768),
	.B1(REGISTERS[423]),
	.B2(FE_OFN12_n2767),
	.ZN(n2245));
   AND4_X1 U2858 (.A1(n2248),
	.A2(n2247),
	.A3(n2246),
	.A4(n2245),
	.ZN(n2265));
   AOI22_X1 U2859 (.A1(REGISTERS[71]),
	.A2(FE_OFN14_n2762),
	.B1(REGISTERS[7]),
	.B2(FE_OFN136_n2761),
	.ZN(n2252));
   AOI22_X1 U2860 (.A1(REGISTERS[199]),
	.A2(FE_OFN55_n2764),
	.B1(REGISTERS[135]),
	.B2(FE_OFN111_n2763),
	.ZN(n2251));
   AOI22_X1 U2861 (.A1(REGISTERS[103]),
	.A2(FE_OFN9_n2766),
	.B1(REGISTERS[39]),
	.B2(FE_OFN52_n2765),
	.ZN(n2250));
   AOI22_X1 U2862 (.A1(REGISTERS[231]),
	.A2(FE_OFN114_n2768),
	.B1(REGISTERS[167]),
	.B2(FE_OFN12_n2767),
	.ZN(n2249));
   AND4_X1 U2863 (.A1(n2252),
	.A2(n2251),
	.A3(n2250),
	.A4(n2249),
	.ZN(n2264));
   AOI22_X1 U2864 (.A1(REGISTERS[839]),
	.A2(FE_OFN14_n2762),
	.B1(REGISTERS[775]),
	.B2(n2761),
	.ZN(n2256));
   AOI22_X1 U2865 (.A1(REGISTERS[967]),
	.A2(FE_OFN56_n2764),
	.B1(REGISTERS[903]),
	.B2(FE_OFN112_n2763),
	.ZN(n2255));
   AOI22_X1 U2866 (.A1(REGISTERS[871]),
	.A2(FE_OFN10_n2766),
	.B1(REGISTERS[807]),
	.B2(FE_OFN53_n2765),
	.ZN(n2254));
   AOI22_X1 U2867 (.A1(REGISTERS[999]),
	.A2(FE_OFN114_n2768),
	.B1(REGISTERS[935]),
	.B2(FE_OFN12_n2767),
	.ZN(n2253));
   NAND4_X1 U2868 (.A1(n2256),
	.A2(n2255),
	.A3(n2254),
	.A4(n2253),
	.ZN(n2262));
   AOI22_X1 U2869 (.A1(REGISTERS[583]),
	.A2(FE_OFN14_n2762),
	.B1(REGISTERS[519]),
	.B2(n2761),
	.ZN(n2260));
   AOI22_X1 U2870 (.A1(REGISTERS[711]),
	.A2(FE_OFN56_n2764),
	.B1(REGISTERS[647]),
	.B2(FE_OFN112_n2763),
	.ZN(n2259));
   AOI22_X1 U2871 (.A1(REGISTERS[615]),
	.A2(FE_OFN10_n2766),
	.B1(REGISTERS[551]),
	.B2(FE_OFN53_n2765),
	.ZN(n2258));
   AOI22_X1 U2872 (.A1(REGISTERS[743]),
	.A2(FE_OFN114_n2768),
	.B1(REGISTERS[679]),
	.B2(FE_OFN12_n2767),
	.ZN(n2257));
   NAND4_X1 U2873 (.A1(n2260),
	.A2(n2259),
	.A3(n2258),
	.A4(n2257),
	.ZN(n2261));
   AOI22_X1 U2874 (.A1(n2262),
	.A2(FE_OFN32_n2776),
	.B1(n2261),
	.B2(FE_OFN30_n2774),
	.ZN(n2263));
   OAI221_X1 U2875 (.A(n2263),
	.B1(n2780),
	.B2(n2265),
	.C1(n2778),
	.C2(n2264),
	.ZN(N55));
   AOI22_X1 U2876 (.A1(REGISTERS[328]),
	.A2(FE_OFN13_n2762),
	.B1(REGISTERS[264]),
	.B2(FE_OFN135_n2761),
	.ZN(n2269));
   AOI22_X1 U2877 (.A1(REGISTERS[456]),
	.A2(n2764),
	.B1(REGISTERS[392]),
	.B2(n2763),
	.ZN(n2268));
   AOI22_X1 U2878 (.A1(REGISTERS[360]),
	.A2(FE_OFN8_n2766),
	.B1(REGISTERS[296]),
	.B2(n2765),
	.ZN(n2267));
   AOI22_X1 U2879 (.A1(REGISTERS[488]),
	.A2(FE_OFN113_n2768),
	.B1(REGISTERS[424]),
	.B2(n2767),
	.ZN(n2266));
   AND4_X1 U2880 (.A1(n2269),
	.A2(n2268),
	.A3(n2267),
	.A4(n2266),
	.ZN(n2286));
   AOI22_X1 U2881 (.A1(REGISTERS[72]),
	.A2(FE_OFN13_n2762),
	.B1(REGISTERS[8]),
	.B2(FE_OFN135_n2761),
	.ZN(n2273));
   AOI22_X1 U2882 (.A1(REGISTERS[200]),
	.A2(n2764),
	.B1(REGISTERS[136]),
	.B2(n2763),
	.ZN(n2272));
   AOI22_X1 U2883 (.A1(REGISTERS[104]),
	.A2(FE_OFN8_n2766),
	.B1(REGISTERS[40]),
	.B2(n2765),
	.ZN(n2271));
   AOI22_X1 U2884 (.A1(REGISTERS[232]),
	.A2(FE_OFN113_n2768),
	.B1(REGISTERS[168]),
	.B2(n2767),
	.ZN(n2270));
   AND4_X1 U2885 (.A1(n2273),
	.A2(n2272),
	.A3(n2271),
	.A4(n2270),
	.ZN(n2285));
   AOI22_X1 U2886 (.A1(REGISTERS[840]),
	.A2(FE_OFN13_n2762),
	.B1(REGISTERS[776]),
	.B2(FE_OFN135_n2761),
	.ZN(n2277));
   AOI22_X1 U2887 (.A1(REGISTERS[968]),
	.A2(FE_OFN54_n2764),
	.B1(REGISTERS[904]),
	.B2(FE_OFN110_n2763),
	.ZN(n2276));
   AOI22_X1 U2888 (.A1(REGISTERS[872]),
	.A2(FE_OFN8_n2766),
	.B1(REGISTERS[808]),
	.B2(n2765),
	.ZN(n2275));
   AOI22_X1 U2889 (.A1(REGISTERS[1000]),
	.A2(n2768),
	.B1(REGISTERS[936]),
	.B2(n2767),
	.ZN(n2274));
   NAND4_X1 U2890 (.A1(n2277),
	.A2(n2276),
	.A3(n2275),
	.A4(n2274),
	.ZN(n2283));
   AOI22_X1 U2891 (.A1(REGISTERS[584]),
	.A2(FE_OFN13_n2762),
	.B1(REGISTERS[520]),
	.B2(FE_OFN135_n2761),
	.ZN(n2281));
   AOI22_X1 U2892 (.A1(REGISTERS[712]),
	.A2(FE_OFN54_n2764),
	.B1(REGISTERS[648]),
	.B2(FE_OFN110_n2763),
	.ZN(n2280));
   AOI22_X1 U2893 (.A1(REGISTERS[616]),
	.A2(FE_OFN8_n2766),
	.B1(REGISTERS[552]),
	.B2(n2765),
	.ZN(n2279));
   AOI22_X1 U2894 (.A1(REGISTERS[744]),
	.A2(n2768),
	.B1(REGISTERS[680]),
	.B2(n2767),
	.ZN(n2278));
   NAND4_X1 U2895 (.A1(n2281),
	.A2(n2280),
	.A3(n2279),
	.A4(n2278),
	.ZN(n2282));
   AOI22_X1 U2896 (.A1(n2283),
	.A2(FE_OFN32_n2776),
	.B1(n2282),
	.B2(FE_OFN30_n2774),
	.ZN(n2284));
   OAI221_X1 U2897 (.A(n2284),
	.B1(n2780),
	.B2(n2286),
	.C1(n2778),
	.C2(n2285),
	.ZN(N54));
   AOI22_X1 U2898 (.A1(REGISTERS[329]),
	.A2(n2762),
	.B1(REGISTERS[265]),
	.B2(n2761),
	.ZN(n2290));
   AOI22_X1 U2899 (.A1(REGISTERS[457]),
	.A2(FE_OFN54_n2764),
	.B1(REGISTERS[393]),
	.B2(FE_OFN110_n2763),
	.ZN(n2289));
   AOI22_X1 U2900 (.A1(REGISTERS[361]),
	.A2(n2766),
	.B1(REGISTERS[297]),
	.B2(n2765),
	.ZN(n2288));
   AOI22_X1 U2901 (.A1(REGISTERS[489]),
	.A2(n2768),
	.B1(REGISTERS[425]),
	.B2(n2767),
	.ZN(n2287));
   AND4_X1 U2902 (.A1(n2290),
	.A2(n2289),
	.A3(n2288),
	.A4(n2287),
	.ZN(n2307));
   AOI22_X1 U2903 (.A1(REGISTERS[73]),
	.A2(n2762),
	.B1(REGISTERS[9]),
	.B2(n2761),
	.ZN(n2294));
   AOI22_X1 U2904 (.A1(REGISTERS[201]),
	.A2(FE_OFN54_n2764),
	.B1(REGISTERS[137]),
	.B2(FE_OFN110_n2763),
	.ZN(n2293));
   AOI22_X1 U2905 (.A1(REGISTERS[105]),
	.A2(n2766),
	.B1(REGISTERS[41]),
	.B2(n2765),
	.ZN(n2292));
   AOI22_X1 U2906 (.A1(REGISTERS[233]),
	.A2(n2768),
	.B1(REGISTERS[169]),
	.B2(n2767),
	.ZN(n2291));
   AND4_X1 U2907 (.A1(n2294),
	.A2(n2293),
	.A3(n2292),
	.A4(n2291),
	.ZN(n2306));
   AOI22_X1 U2908 (.A1(REGISTERS[841]),
	.A2(n2762),
	.B1(REGISTERS[777]),
	.B2(n2761),
	.ZN(n2298));
   AOI22_X1 U2909 (.A1(REGISTERS[969]),
	.A2(FE_OFN54_n2764),
	.B1(REGISTERS[905]),
	.B2(n2763),
	.ZN(n2297));
   AOI22_X1 U2910 (.A1(REGISTERS[873]),
	.A2(FE_OFN9_n2766),
	.B1(REGISTERS[809]),
	.B2(FE_OFN53_n2765),
	.ZN(n2296));
   AOI22_X1 U2911 (.A1(REGISTERS[1001]),
	.A2(n2768),
	.B1(REGISTERS[937]),
	.B2(n2767),
	.ZN(n2295));
   NAND4_X1 U2912 (.A1(n2298),
	.A2(n2297),
	.A3(n2296),
	.A4(n2295),
	.ZN(n2304));
   AOI22_X1 U2913 (.A1(REGISTERS[585]),
	.A2(n2762),
	.B1(REGISTERS[521]),
	.B2(n2761),
	.ZN(n2302));
   AOI22_X1 U2914 (.A1(REGISTERS[713]),
	.A2(FE_OFN54_n2764),
	.B1(REGISTERS[649]),
	.B2(n2763),
	.ZN(n2301));
   AOI22_X1 U2915 (.A1(REGISTERS[617]),
	.A2(FE_OFN9_n2766),
	.B1(REGISTERS[553]),
	.B2(FE_OFN53_n2765),
	.ZN(n2300));
   AOI22_X1 U2916 (.A1(REGISTERS[745]),
	.A2(n2768),
	.B1(REGISTERS[681]),
	.B2(n2767),
	.ZN(n2299));
   NAND4_X1 U2917 (.A1(n2302),
	.A2(n2301),
	.A3(n2300),
	.A4(n2299),
	.ZN(n2303));
   AOI22_X1 U2918 (.A1(n2304),
	.A2(FE_OFN32_n2776),
	.B1(n2303),
	.B2(FE_OFN30_n2774),
	.ZN(n2305));
   OAI221_X1 U2919 (.A(n2305),
	.B1(n2780),
	.B2(n2307),
	.C1(n2778),
	.C2(n2306),
	.ZN(N53));
   AOI22_X1 U2920 (.A1(REGISTERS[330]),
	.A2(n2762),
	.B1(REGISTERS[266]),
	.B2(FE_OFN135_n2761),
	.ZN(n2311));
   AOI22_X1 U2921 (.A1(REGISTERS[458]),
	.A2(n2764),
	.B1(REGISTERS[394]),
	.B2(n2763),
	.ZN(n2310));
   AOI22_X1 U2922 (.A1(REGISTERS[362]),
	.A2(FE_OFN8_n2766),
	.B1(REGISTERS[298]),
	.B2(n2765),
	.ZN(n2309));
   AOI22_X1 U2923 (.A1(REGISTERS[490]),
	.A2(n2768),
	.B1(REGISTERS[426]),
	.B2(n2767),
	.ZN(n2308));
   AND4_X1 U2924 (.A1(n2311),
	.A2(n2310),
	.A3(n2309),
	.A4(n2308),
	.ZN(n2328));
   AOI22_X1 U2925 (.A1(REGISTERS[74]),
	.A2(n2762),
	.B1(REGISTERS[10]),
	.B2(n2761),
	.ZN(n2315));
   AOI22_X1 U2926 (.A1(REGISTERS[202]),
	.A2(n2764),
	.B1(REGISTERS[138]),
	.B2(n2763),
	.ZN(n2314));
   AOI22_X1 U2927 (.A1(REGISTERS[106]),
	.A2(FE_OFN8_n2766),
	.B1(REGISTERS[42]),
	.B2(n2765),
	.ZN(n2313));
   AOI22_X1 U2928 (.A1(REGISTERS[234]),
	.A2(n2768),
	.B1(REGISTERS[170]),
	.B2(n2767),
	.ZN(n2312));
   AND4_X1 U2929 (.A1(n2315),
	.A2(n2314),
	.A3(n2313),
	.A4(n2312),
	.ZN(n2327));
   AOI22_X1 U2930 (.A1(REGISTERS[842]),
	.A2(n2762),
	.B1(REGISTERS[778]),
	.B2(n2761),
	.ZN(n2319));
   AOI22_X1 U2931 (.A1(REGISTERS[970]),
	.A2(FE_OFN54_n2764),
	.B1(REGISTERS[906]),
	.B2(FE_OFN110_n2763),
	.ZN(n2318));
   AOI22_X1 U2932 (.A1(REGISTERS[874]),
	.A2(n2766),
	.B1(REGISTERS[810]),
	.B2(n2765),
	.ZN(n2317));
   AOI22_X1 U2933 (.A1(REGISTERS[1002]),
	.A2(n2768),
	.B1(REGISTERS[938]),
	.B2(n2767),
	.ZN(n2316));
   NAND4_X1 U2934 (.A1(n2319),
	.A2(n2318),
	.A3(n2317),
	.A4(n2316),
	.ZN(n2325));
   AOI22_X1 U2935 (.A1(REGISTERS[586]),
	.A2(n2762),
	.B1(REGISTERS[522]),
	.B2(n2761),
	.ZN(n2323));
   AOI22_X1 U2936 (.A1(REGISTERS[714]),
	.A2(FE_OFN54_n2764),
	.B1(REGISTERS[650]),
	.B2(FE_OFN110_n2763),
	.ZN(n2322));
   AOI22_X1 U2937 (.A1(REGISTERS[618]),
	.A2(n2766),
	.B1(REGISTERS[554]),
	.B2(n2765),
	.ZN(n2321));
   AOI22_X1 U2938 (.A1(REGISTERS[746]),
	.A2(n2768),
	.B1(REGISTERS[682]),
	.B2(n2767),
	.ZN(n2320));
   NAND4_X1 U2939 (.A1(n2323),
	.A2(n2322),
	.A3(n2321),
	.A4(n2320),
	.ZN(n2324));
   AOI22_X1 U2940 (.A1(n2325),
	.A2(FE_OFN32_n2776),
	.B1(n2324),
	.B2(FE_OFN30_n2774),
	.ZN(n2326));
   OAI221_X1 U2941 (.A(n2326),
	.B1(n2780),
	.B2(n2328),
	.C1(n2778),
	.C2(n2327),
	.ZN(N52));
   AOI22_X1 U2942 (.A1(REGISTERS[331]),
	.A2(n2762),
	.B1(REGISTERS[267]),
	.B2(n2761),
	.ZN(n2332));
   AOI22_X1 U2943 (.A1(REGISTERS[459]),
	.A2(FE_OFN54_n2764),
	.B1(REGISTERS[395]),
	.B2(n2763),
	.ZN(n2331));
   AOI22_X1 U2944 (.A1(REGISTERS[363]),
	.A2(FE_OFN9_n2766),
	.B1(REGISTERS[299]),
	.B2(FE_OFN53_n2765),
	.ZN(n2330));
   AOI22_X1 U2945 (.A1(REGISTERS[491]),
	.A2(n2768),
	.B1(REGISTERS[427]),
	.B2(n2767),
	.ZN(n2329));
   AND4_X1 U2946 (.A1(n2332),
	.A2(n2331),
	.A3(n2330),
	.A4(n2329),
	.ZN(n2349));
   AOI22_X1 U2947 (.A1(REGISTERS[75]),
	.A2(n2762),
	.B1(REGISTERS[11]),
	.B2(n2761),
	.ZN(n2336));
   AOI22_X1 U2948 (.A1(REGISTERS[203]),
	.A2(FE_OFN54_n2764),
	.B1(REGISTERS[139]),
	.B2(n2763),
	.ZN(n2335));
   AOI22_X1 U2949 (.A1(REGISTERS[107]),
	.A2(FE_OFN9_n2766),
	.B1(REGISTERS[43]),
	.B2(FE_OFN53_n2765),
	.ZN(n2334));
   AOI22_X1 U2950 (.A1(REGISTERS[235]),
	.A2(n2768),
	.B1(REGISTERS[171]),
	.B2(n2767),
	.ZN(n2333));
   AND4_X1 U2951 (.A1(n2336),
	.A2(n2335),
	.A3(n2334),
	.A4(n2333),
	.ZN(n2348));
   AOI22_X1 U2952 (.A1(REGISTERS[843]),
	.A2(n2762),
	.B1(REGISTERS[779]),
	.B2(n2761),
	.ZN(n2340));
   AOI22_X1 U2953 (.A1(REGISTERS[971]),
	.A2(FE_OFN54_n2764),
	.B1(REGISTERS[907]),
	.B2(n2763),
	.ZN(n2339));
   AOI22_X1 U2954 (.A1(REGISTERS[875]),
	.A2(FE_OFN9_n2766),
	.B1(REGISTERS[811]),
	.B2(FE_OFN53_n2765),
	.ZN(n2338));
   AOI22_X1 U2955 (.A1(REGISTERS[1003]),
	.A2(n2768),
	.B1(REGISTERS[939]),
	.B2(n2767),
	.ZN(n2337));
   NAND4_X1 U2956 (.A1(n2340),
	.A2(n2339),
	.A3(n2338),
	.A4(n2337),
	.ZN(n2346));
   AOI22_X1 U2957 (.A1(REGISTERS[587]),
	.A2(n2762),
	.B1(REGISTERS[523]),
	.B2(n2761),
	.ZN(n2344));
   AOI22_X1 U2958 (.A1(REGISTERS[715]),
	.A2(FE_OFN54_n2764),
	.B1(REGISTERS[651]),
	.B2(n2763),
	.ZN(n2343));
   AOI22_X1 U2959 (.A1(REGISTERS[619]),
	.A2(FE_OFN9_n2766),
	.B1(REGISTERS[555]),
	.B2(FE_OFN53_n2765),
	.ZN(n2342));
   AOI22_X1 U2960 (.A1(REGISTERS[747]),
	.A2(n2768),
	.B1(REGISTERS[683]),
	.B2(n2767),
	.ZN(n2341));
   NAND4_X1 U2961 (.A1(n2344),
	.A2(n2343),
	.A3(n2342),
	.A4(n2341),
	.ZN(n2345));
   AOI22_X1 U2962 (.A1(n2346),
	.A2(FE_OFN32_n2776),
	.B1(n2345),
	.B2(FE_OFN30_n2774),
	.ZN(n2347));
   OAI221_X1 U2963 (.A(n2347),
	.B1(n2780),
	.B2(n2349),
	.C1(n2778),
	.C2(n2348),
	.ZN(N51));
   AOI22_X1 U2964 (.A1(REGISTERS[332]),
	.A2(n2762),
	.B1(REGISTERS[268]),
	.B2(n2761),
	.ZN(n2353));
   AOI22_X1 U2965 (.A1(REGISTERS[460]),
	.A2(n2764),
	.B1(REGISTERS[396]),
	.B2(n2763),
	.ZN(n2352));
   AOI22_X1 U2966 (.A1(REGISTERS[364]),
	.A2(FE_OFN8_n2766),
	.B1(REGISTERS[300]),
	.B2(n2765),
	.ZN(n2351));
   AOI22_X1 U2967 (.A1(REGISTERS[492]),
	.A2(n2768),
	.B1(REGISTERS[428]),
	.B2(n2767),
	.ZN(n2350));
   AND4_X1 U2968 (.A1(n2353),
	.A2(n2352),
	.A3(n2351),
	.A4(n2350),
	.ZN(n2370));
   AOI22_X1 U2969 (.A1(REGISTERS[76]),
	.A2(n2762),
	.B1(REGISTERS[12]),
	.B2(n2761),
	.ZN(n2357));
   AOI22_X1 U2970 (.A1(REGISTERS[204]),
	.A2(n2764),
	.B1(REGISTERS[140]),
	.B2(n2763),
	.ZN(n2356));
   AOI22_X1 U2971 (.A1(REGISTERS[108]),
	.A2(FE_OFN8_n2766),
	.B1(REGISTERS[44]),
	.B2(n2765),
	.ZN(n2355));
   AOI22_X1 U2972 (.A1(REGISTERS[236]),
	.A2(n2768),
	.B1(REGISTERS[172]),
	.B2(n2767),
	.ZN(n2354));
   AND4_X1 U2973 (.A1(n2357),
	.A2(n2356),
	.A3(n2355),
	.A4(n2354),
	.ZN(n2369));
   AOI22_X1 U2974 (.A1(REGISTERS[844]),
	.A2(n2762),
	.B1(REGISTERS[780]),
	.B2(n2761),
	.ZN(n2361));
   AOI22_X1 U2975 (.A1(REGISTERS[972]),
	.A2(FE_OFN54_n2764),
	.B1(REGISTERS[908]),
	.B2(FE_OFN110_n2763),
	.ZN(n2360));
   AOI22_X1 U2976 (.A1(REGISTERS[876]),
	.A2(n2766),
	.B1(REGISTERS[812]),
	.B2(n2765),
	.ZN(n2359));
   AOI22_X1 U2977 (.A1(REGISTERS[1004]),
	.A2(n2768),
	.B1(REGISTERS[940]),
	.B2(n2767),
	.ZN(n2358));
   NAND4_X1 U2978 (.A1(n2361),
	.A2(n2360),
	.A3(n2359),
	.A4(n2358),
	.ZN(n2367));
   AOI22_X1 U2979 (.A1(REGISTERS[588]),
	.A2(n2762),
	.B1(REGISTERS[524]),
	.B2(n2761),
	.ZN(n2365));
   AOI22_X1 U2980 (.A1(REGISTERS[716]),
	.A2(FE_OFN54_n2764),
	.B1(REGISTERS[652]),
	.B2(FE_OFN110_n2763),
	.ZN(n2364));
   AOI22_X1 U2981 (.A1(REGISTERS[620]),
	.A2(n2766),
	.B1(REGISTERS[556]),
	.B2(n2765),
	.ZN(n2363));
   AOI22_X1 U2982 (.A1(REGISTERS[748]),
	.A2(n2768),
	.B1(REGISTERS[684]),
	.B2(n2767),
	.ZN(n2362));
   NAND4_X1 U2983 (.A1(n2365),
	.A2(n2364),
	.A3(n2363),
	.A4(n2362),
	.ZN(n2366));
   AOI22_X1 U2984 (.A1(n2367),
	.A2(FE_OFN32_n2776),
	.B1(n2366),
	.B2(FE_OFN30_n2774),
	.ZN(n2368));
   OAI221_X1 U2985 (.A(n2368),
	.B1(n2780),
	.B2(n2370),
	.C1(n2778),
	.C2(n2369),
	.ZN(N50));
   AOI22_X1 U2986 (.A1(REGISTERS[333]),
	.A2(FE_OFN13_n2762),
	.B1(REGISTERS[269]),
	.B2(FE_OFN135_n2761),
	.ZN(n2374));
   AOI22_X1 U2987 (.A1(REGISTERS[461]),
	.A2(n2764),
	.B1(REGISTERS[397]),
	.B2(n2763),
	.ZN(n2373));
   AOI22_X1 U2988 (.A1(REGISTERS[365]),
	.A2(FE_OFN8_n2766),
	.B1(REGISTERS[301]),
	.B2(FE_OFN51_n2765),
	.ZN(n2372));
   AOI22_X1 U2989 (.A1(REGISTERS[493]),
	.A2(FE_OFN113_n2768),
	.B1(REGISTERS[429]),
	.B2(n2767),
	.ZN(n2371));
   AND4_X1 U2990 (.A1(n2374),
	.A2(n2373),
	.A3(n2372),
	.A4(n2371),
	.ZN(n2391));
   AOI22_X1 U2991 (.A1(REGISTERS[77]),
	.A2(FE_OFN13_n2762),
	.B1(REGISTERS[13]),
	.B2(FE_OFN135_n2761),
	.ZN(n2378));
   AOI22_X1 U2992 (.A1(REGISTERS[205]),
	.A2(n2764),
	.B1(REGISTERS[141]),
	.B2(n2763),
	.ZN(n2377));
   AOI22_X1 U2993 (.A1(REGISTERS[109]),
	.A2(FE_OFN8_n2766),
	.B1(REGISTERS[45]),
	.B2(FE_OFN51_n2765),
	.ZN(n2376));
   AOI22_X1 U2994 (.A1(REGISTERS[237]),
	.A2(FE_OFN113_n2768),
	.B1(REGISTERS[173]),
	.B2(FE_OFN11_n2767),
	.ZN(n2375));
   AND4_X1 U2995 (.A1(n2378),
	.A2(n2377),
	.A3(n2376),
	.A4(n2375),
	.ZN(n2390));
   AOI22_X1 U2996 (.A1(REGISTERS[845]),
	.A2(FE_OFN13_n2762),
	.B1(REGISTERS[781]),
	.B2(FE_OFN135_n2761),
	.ZN(n2382));
   AOI22_X1 U2997 (.A1(REGISTERS[973]),
	.A2(FE_OFN54_n2764),
	.B1(REGISTERS[909]),
	.B2(FE_OFN110_n2763),
	.ZN(n2381));
   AOI22_X1 U2998 (.A1(REGISTERS[877]),
	.A2(FE_OFN8_n2766),
	.B1(REGISTERS[813]),
	.B2(n2765),
	.ZN(n2380));
   AOI22_X1 U2999 (.A1(REGISTERS[1005]),
	.A2(FE_OFN113_n2768),
	.B1(REGISTERS[941]),
	.B2(FE_OFN11_n2767),
	.ZN(n2379));
   NAND4_X1 U3000 (.A1(n2382),
	.A2(n2381),
	.A3(n2380),
	.A4(n2379),
	.ZN(n2388));
   AOI22_X1 U3001 (.A1(REGISTERS[589]),
	.A2(FE_OFN13_n2762),
	.B1(REGISTERS[525]),
	.B2(FE_OFN135_n2761),
	.ZN(n2386));
   AOI22_X1 U3002 (.A1(REGISTERS[717]),
	.A2(FE_OFN54_n2764),
	.B1(REGISTERS[653]),
	.B2(FE_OFN110_n2763),
	.ZN(n2385));
   AOI22_X1 U3003 (.A1(REGISTERS[621]),
	.A2(FE_OFN9_n2766),
	.B1(REGISTERS[557]),
	.B2(n2765),
	.ZN(n2384));
   AOI22_X1 U3004 (.A1(REGISTERS[749]),
	.A2(FE_OFN113_n2768),
	.B1(REGISTERS[685]),
	.B2(FE_OFN11_n2767),
	.ZN(n2383));
   NAND4_X1 U3005 (.A1(n2386),
	.A2(n2385),
	.A3(n2384),
	.A4(n2383),
	.ZN(n2387));
   AOI22_X1 U3006 (.A1(n2388),
	.A2(FE_OFN32_n2776),
	.B1(n2387),
	.B2(FE_OFN30_n2774),
	.ZN(n2389));
   OAI221_X1 U3007 (.A(n2389),
	.B1(n2780),
	.B2(n2391),
	.C1(n2778),
	.C2(n2390),
	.ZN(N49));
   AOI22_X1 U3008 (.A1(REGISTERS[334]),
	.A2(FE_OFN14_n2762),
	.B1(REGISTERS[270]),
	.B2(FE_OFN136_n2761),
	.ZN(n2395));
   AOI22_X1 U3009 (.A1(REGISTERS[462]),
	.A2(FE_OFN54_n2764),
	.B1(REGISTERS[398]),
	.B2(FE_OFN111_n2763),
	.ZN(n2394));
   AOI22_X1 U3010 (.A1(REGISTERS[366]),
	.A2(FE_OFN9_n2766),
	.B1(REGISTERS[302]),
	.B2(FE_OFN53_n2765),
	.ZN(n2393));
   AOI22_X1 U3011 (.A1(REGISTERS[494]),
	.A2(FE_OFN114_n2768),
	.B1(REGISTERS[430]),
	.B2(FE_OFN12_n2767),
	.ZN(n2392));
   AND4_X1 U3012 (.A1(n2395),
	.A2(n2394),
	.A3(n2393),
	.A4(n2392),
	.ZN(n2412));
   AOI22_X1 U3013 (.A1(REGISTERS[78]),
	.A2(FE_OFN14_n2762),
	.B1(REGISTERS[14]),
	.B2(FE_OFN136_n2761),
	.ZN(n2399));
   AOI22_X1 U3014 (.A1(REGISTERS[206]),
	.A2(FE_OFN54_n2764),
	.B1(REGISTERS[142]),
	.B2(FE_OFN111_n2763),
	.ZN(n2398));
   AOI22_X1 U3015 (.A1(REGISTERS[110]),
	.A2(FE_OFN9_n2766),
	.B1(REGISTERS[46]),
	.B2(FE_OFN53_n2765),
	.ZN(n2397));
   AOI22_X1 U3016 (.A1(REGISTERS[238]),
	.A2(FE_OFN114_n2768),
	.B1(REGISTERS[174]),
	.B2(FE_OFN12_n2767),
	.ZN(n2396));
   AND4_X1 U3017 (.A1(n2399),
	.A2(n2398),
	.A3(n2397),
	.A4(n2396),
	.ZN(n2411));
   AOI22_X1 U3018 (.A1(REGISTERS[846]),
	.A2(FE_OFN14_n2762),
	.B1(REGISTERS[782]),
	.B2(n2761),
	.ZN(n2403));
   AOI22_X1 U3019 (.A1(REGISTERS[974]),
	.A2(FE_OFN56_n2764),
	.B1(REGISTERS[910]),
	.B2(FE_OFN112_n2763),
	.ZN(n2402));
   AOI22_X1 U3020 (.A1(REGISTERS[878]),
	.A2(FE_OFN9_n2766),
	.B1(REGISTERS[814]),
	.B2(FE_OFN53_n2765),
	.ZN(n2401));
   AOI22_X1 U3021 (.A1(REGISTERS[1006]),
	.A2(FE_OFN114_n2768),
	.B1(REGISTERS[942]),
	.B2(FE_OFN12_n2767),
	.ZN(n2400));
   NAND4_X1 U3022 (.A1(n2403),
	.A2(n2402),
	.A3(n2401),
	.A4(n2400),
	.ZN(n2409));
   AOI22_X1 U3023 (.A1(REGISTERS[590]),
	.A2(FE_OFN14_n2762),
	.B1(REGISTERS[526]),
	.B2(n2761),
	.ZN(n2407));
   AOI22_X1 U3024 (.A1(REGISTERS[718]),
	.A2(FE_OFN56_n2764),
	.B1(REGISTERS[654]),
	.B2(FE_OFN112_n2763),
	.ZN(n2406));
   AOI22_X1 U3025 (.A1(REGISTERS[622]),
	.A2(FE_OFN9_n2766),
	.B1(REGISTERS[558]),
	.B2(FE_OFN53_n2765),
	.ZN(n2405));
   AOI22_X1 U3026 (.A1(REGISTERS[750]),
	.A2(FE_OFN114_n2768),
	.B1(REGISTERS[686]),
	.B2(FE_OFN12_n2767),
	.ZN(n2404));
   NAND4_X1 U3027 (.A1(n2407),
	.A2(n2406),
	.A3(n2405),
	.A4(n2404),
	.ZN(n2408));
   AOI22_X1 U3028 (.A1(n2409),
	.A2(FE_OFN32_n2776),
	.B1(n2408),
	.B2(FE_OFN30_n2774),
	.ZN(n2410));
   OAI221_X1 U3029 (.A(n2410),
	.B1(n2780),
	.B2(n2412),
	.C1(n2778),
	.C2(n2411),
	.ZN(N48));
   AOI22_X1 U3030 (.A1(REGISTERS[335]),
	.A2(n2762),
	.B1(REGISTERS[271]),
	.B2(n2761),
	.ZN(n2416));
   AOI22_X1 U3031 (.A1(REGISTERS[463]),
	.A2(n2764),
	.B1(REGISTERS[399]),
	.B2(n2763),
	.ZN(n2415));
   AOI22_X1 U3032 (.A1(REGISTERS[367]),
	.A2(n2766),
	.B1(REGISTERS[303]),
	.B2(n2765),
	.ZN(n2414));
   AOI22_X1 U3033 (.A1(REGISTERS[495]),
	.A2(n2768),
	.B1(REGISTERS[431]),
	.B2(n2767),
	.ZN(n2413));
   AND4_X1 U3034 (.A1(n2416),
	.A2(n2415),
	.A3(n2414),
	.A4(n2413),
	.ZN(n2433));
   AOI22_X1 U3035 (.A1(REGISTERS[79]),
	.A2(n2762),
	.B1(REGISTERS[15]),
	.B2(n2761),
	.ZN(n2420));
   AOI22_X1 U3036 (.A1(REGISTERS[207]),
	.A2(n2764),
	.B1(REGISTERS[143]),
	.B2(n2763),
	.ZN(n2419));
   AOI22_X1 U3037 (.A1(REGISTERS[111]),
	.A2(FE_OFN8_n2766),
	.B1(REGISTERS[47]),
	.B2(n2765),
	.ZN(n2418));
   AOI22_X1 U3038 (.A1(REGISTERS[239]),
	.A2(n2768),
	.B1(REGISTERS[175]),
	.B2(n2767),
	.ZN(n2417));
   AND4_X1 U3039 (.A1(n2420),
	.A2(n2419),
	.A3(n2418),
	.A4(n2417),
	.ZN(n2432));
   AOI22_X1 U3040 (.A1(REGISTERS[847]),
	.A2(n2762),
	.B1(REGISTERS[783]),
	.B2(n2761),
	.ZN(n2424));
   AOI22_X1 U3041 (.A1(REGISTERS[975]),
	.A2(FE_OFN56_n2764),
	.B1(REGISTERS[911]),
	.B2(FE_OFN112_n2763),
	.ZN(n2423));
   AOI22_X1 U3042 (.A1(REGISTERS[879]),
	.A2(FE_OFN9_n2766),
	.B1(REGISTERS[815]),
	.B2(FE_OFN53_n2765),
	.ZN(n2422));
   AOI22_X1 U3043 (.A1(REGISTERS[1007]),
	.A2(FE_OFN114_n2768),
	.B1(REGISTERS[943]),
	.B2(FE_OFN12_n2767),
	.ZN(n2421));
   NAND4_X1 U3044 (.A1(n2424),
	.A2(n2423),
	.A3(n2422),
	.A4(n2421),
	.ZN(n2430));
   AOI22_X1 U3045 (.A1(REGISTERS[591]),
	.A2(n2762),
	.B1(REGISTERS[527]),
	.B2(n2761),
	.ZN(n2428));
   AOI22_X1 U3046 (.A1(REGISTERS[719]),
	.A2(FE_OFN56_n2764),
	.B1(REGISTERS[655]),
	.B2(FE_OFN112_n2763),
	.ZN(n2427));
   AOI22_X1 U3047 (.A1(REGISTERS[623]),
	.A2(FE_OFN9_n2766),
	.B1(REGISTERS[559]),
	.B2(FE_OFN53_n2765),
	.ZN(n2426));
   AOI22_X1 U3048 (.A1(REGISTERS[751]),
	.A2(FE_OFN114_n2768),
	.B1(REGISTERS[687]),
	.B2(FE_OFN12_n2767),
	.ZN(n2425));
   NAND4_X1 U3049 (.A1(n2428),
	.A2(n2427),
	.A3(n2426),
	.A4(n2425),
	.ZN(n2429));
   AOI22_X1 U3050 (.A1(n2430),
	.A2(FE_OFN32_n2776),
	.B1(n2429),
	.B2(FE_OFN30_n2774),
	.ZN(n2431));
   OAI221_X1 U3051 (.A(n2431),
	.B1(n2780),
	.B2(n2433),
	.C1(n2778),
	.C2(n2432),
	.ZN(N47));
   AOI22_X1 U3052 (.A1(REGISTERS[336]),
	.A2(n2762),
	.B1(REGISTERS[272]),
	.B2(n2761),
	.ZN(n2437));
   AOI22_X1 U3053 (.A1(REGISTERS[464]),
	.A2(FE_OFN54_n2764),
	.B1(REGISTERS[400]),
	.B2(n2763),
	.ZN(n2436));
   AOI22_X1 U3054 (.A1(REGISTERS[368]),
	.A2(FE_OFN9_n2766),
	.B1(REGISTERS[304]),
	.B2(FE_OFN53_n2765),
	.ZN(n2435));
   AOI22_X1 U3055 (.A1(REGISTERS[496]),
	.A2(n2768),
	.B1(REGISTERS[432]),
	.B2(n2767),
	.ZN(n2434));
   AND4_X1 U3056 (.A1(n2437),
	.A2(n2436),
	.A3(n2435),
	.A4(n2434),
	.ZN(n2454));
   AOI22_X1 U3057 (.A1(REGISTERS[80]),
	.A2(n2762),
	.B1(REGISTERS[16]),
	.B2(n2761),
	.ZN(n2441));
   AOI22_X1 U3058 (.A1(REGISTERS[208]),
	.A2(FE_OFN54_n2764),
	.B1(REGISTERS[144]),
	.B2(n2763),
	.ZN(n2440));
   AOI22_X1 U3059 (.A1(REGISTERS[112]),
	.A2(FE_OFN9_n2766),
	.B1(REGISTERS[48]),
	.B2(FE_OFN53_n2765),
	.ZN(n2439));
   AOI22_X1 U3060 (.A1(REGISTERS[240]),
	.A2(n2768),
	.B1(REGISTERS[176]),
	.B2(n2767),
	.ZN(n2438));
   AND4_X1 U3061 (.A1(n2441),
	.A2(n2440),
	.A3(n2439),
	.A4(n2438),
	.ZN(n2453));
   AOI22_X1 U3062 (.A1(REGISTERS[848]),
	.A2(n2762),
	.B1(REGISTERS[784]),
	.B2(n2761),
	.ZN(n2445));
   AOI22_X1 U3063 (.A1(REGISTERS[976]),
	.A2(FE_OFN56_n2764),
	.B1(REGISTERS[912]),
	.B2(FE_OFN112_n2763),
	.ZN(n2444));
   AOI22_X1 U3064 (.A1(REGISTERS[880]),
	.A2(FE_OFN9_n2766),
	.B1(REGISTERS[816]),
	.B2(FE_OFN53_n2765),
	.ZN(n2443));
   AOI22_X1 U3065 (.A1(REGISTERS[1008]),
	.A2(FE_OFN114_n2768),
	.B1(REGISTERS[944]),
	.B2(FE_OFN12_n2767),
	.ZN(n2442));
   NAND4_X1 U3066 (.A1(n2445),
	.A2(n2444),
	.A3(n2443),
	.A4(n2442),
	.ZN(n2451));
   AOI22_X1 U3067 (.A1(REGISTERS[592]),
	.A2(n2762),
	.B1(REGISTERS[528]),
	.B2(n2761),
	.ZN(n2449));
   AOI22_X1 U3068 (.A1(REGISTERS[720]),
	.A2(FE_OFN54_n2764),
	.B1(REGISTERS[656]),
	.B2(n2763),
	.ZN(n2448));
   AOI22_X1 U3069 (.A1(REGISTERS[624]),
	.A2(FE_OFN9_n2766),
	.B1(REGISTERS[560]),
	.B2(FE_OFN53_n2765),
	.ZN(n2447));
   AOI22_X1 U3070 (.A1(REGISTERS[752]),
	.A2(n2768),
	.B1(REGISTERS[688]),
	.B2(FE_OFN12_n2767),
	.ZN(n2446));
   NAND4_X1 U3071 (.A1(n2449),
	.A2(n2448),
	.A3(n2447),
	.A4(n2446),
	.ZN(n2450));
   AOI22_X1 U3072 (.A1(n2451),
	.A2(FE_OFN32_n2776),
	.B1(n2450),
	.B2(FE_OFN30_n2774),
	.ZN(n2452));
   OAI221_X1 U3073 (.A(n2452),
	.B1(n2780),
	.B2(n2454),
	.C1(n2778),
	.C2(n2453),
	.ZN(N46));
   AOI22_X1 U3074 (.A1(REGISTERS[337]),
	.A2(FE_OFN14_n2762),
	.B1(REGISTERS[273]),
	.B2(FE_OFN136_n2761),
	.ZN(n2458));
   AOI22_X1 U3075 (.A1(REGISTERS[465]),
	.A2(FE_OFN55_n2764),
	.B1(REGISTERS[401]),
	.B2(FE_OFN111_n2763),
	.ZN(n2457));
   AOI22_X1 U3076 (.A1(REGISTERS[369]),
	.A2(FE_OFN9_n2766),
	.B1(REGISTERS[305]),
	.B2(FE_OFN52_n2765),
	.ZN(n2456));
   AOI22_X1 U3077 (.A1(REGISTERS[497]),
	.A2(FE_OFN114_n2768),
	.B1(REGISTERS[433]),
	.B2(FE_OFN12_n2767),
	.ZN(n2455));
   AND4_X1 U3078 (.A1(n2458),
	.A2(n2457),
	.A3(n2456),
	.A4(n2455),
	.ZN(n2475));
   AOI22_X1 U3079 (.A1(REGISTERS[81]),
	.A2(FE_OFN14_n2762),
	.B1(REGISTERS[17]),
	.B2(FE_OFN136_n2761),
	.ZN(n2462));
   AOI22_X1 U3080 (.A1(REGISTERS[209]),
	.A2(FE_OFN55_n2764),
	.B1(REGISTERS[145]),
	.B2(FE_OFN111_n2763),
	.ZN(n2461));
   AOI22_X1 U3081 (.A1(REGISTERS[113]),
	.A2(FE_OFN9_n2766),
	.B1(REGISTERS[49]),
	.B2(FE_OFN52_n2765),
	.ZN(n2460));
   AOI22_X1 U3082 (.A1(REGISTERS[241]),
	.A2(FE_OFN114_n2768),
	.B1(REGISTERS[177]),
	.B2(FE_OFN12_n2767),
	.ZN(n2459));
   AND4_X1 U3083 (.A1(n2462),
	.A2(n2461),
	.A3(n2460),
	.A4(n2459),
	.ZN(n2474));
   AOI22_X1 U3084 (.A1(REGISTERS[849]),
	.A2(FE_OFN14_n2762),
	.B1(REGISTERS[785]),
	.B2(FE_OFN136_n2761),
	.ZN(n2466));
   AOI22_X1 U3085 (.A1(REGISTERS[977]),
	.A2(FE_OFN56_n2764),
	.B1(REGISTERS[913]),
	.B2(FE_OFN112_n2763),
	.ZN(n2465));
   AOI22_X1 U3086 (.A1(REGISTERS[881]),
	.A2(FE_OFN10_n2766),
	.B1(REGISTERS[817]),
	.B2(FE_OFN53_n2765),
	.ZN(n2464));
   AOI22_X1 U3087 (.A1(REGISTERS[1009]),
	.A2(FE_OFN114_n2768),
	.B1(REGISTERS[945]),
	.B2(FE_OFN12_n2767),
	.ZN(n2463));
   NAND4_X1 U3088 (.A1(n2466),
	.A2(n2465),
	.A3(n2464),
	.A4(n2463),
	.ZN(n2472));
   AOI22_X1 U3089 (.A1(REGISTERS[593]),
	.A2(FE_OFN14_n2762),
	.B1(REGISTERS[529]),
	.B2(FE_OFN136_n2761),
	.ZN(n2470));
   AOI22_X1 U3090 (.A1(REGISTERS[721]),
	.A2(FE_OFN56_n2764),
	.B1(REGISTERS[657]),
	.B2(FE_OFN112_n2763),
	.ZN(n2469));
   AOI22_X1 U3091 (.A1(REGISTERS[625]),
	.A2(FE_OFN10_n2766),
	.B1(REGISTERS[561]),
	.B2(FE_OFN53_n2765),
	.ZN(n2468));
   AOI22_X1 U3092 (.A1(REGISTERS[753]),
	.A2(FE_OFN114_n2768),
	.B1(REGISTERS[689]),
	.B2(FE_OFN12_n2767),
	.ZN(n2467));
   NAND4_X1 U3093 (.A1(n2470),
	.A2(n2469),
	.A3(n2468),
	.A4(n2467),
	.ZN(n2471));
   AOI22_X1 U3094 (.A1(n2472),
	.A2(FE_OFN32_n2776),
	.B1(n2471),
	.B2(FE_OFN30_n2774),
	.ZN(n2473));
   OAI221_X1 U3095 (.A(n2473),
	.B1(n2780),
	.B2(n2475),
	.C1(n2778),
	.C2(n2474),
	.ZN(N45));
   AOI22_X1 U3096 (.A1(REGISTERS[338]),
	.A2(FE_OFN13_n2762),
	.B1(REGISTERS[274]),
	.B2(FE_OFN135_n2761),
	.ZN(n2479));
   AOI22_X1 U3097 (.A1(REGISTERS[466]),
	.A2(n2764),
	.B1(REGISTERS[402]),
	.B2(n2763),
	.ZN(n2478));
   AOI22_X1 U3098 (.A1(REGISTERS[370]),
	.A2(FE_OFN8_n2766),
	.B1(REGISTERS[306]),
	.B2(FE_OFN51_n2765),
	.ZN(n2477));
   AOI22_X1 U3099 (.A1(REGISTERS[498]),
	.A2(FE_OFN113_n2768),
	.B1(REGISTERS[434]),
	.B2(FE_OFN11_n2767),
	.ZN(n2476));
   AND4_X1 U3100 (.A1(n2479),
	.A2(n2478),
	.A3(n2477),
	.A4(n2476),
	.ZN(n2496));
   AOI22_X1 U3101 (.A1(REGISTERS[82]),
	.A2(FE_OFN13_n2762),
	.B1(REGISTERS[18]),
	.B2(FE_OFN135_n2761),
	.ZN(n2483));
   AOI22_X1 U3102 (.A1(REGISTERS[210]),
	.A2(n2764),
	.B1(REGISTERS[146]),
	.B2(n2763),
	.ZN(n2482));
   AOI22_X1 U3103 (.A1(REGISTERS[114]),
	.A2(FE_OFN8_n2766),
	.B1(REGISTERS[50]),
	.B2(FE_OFN51_n2765),
	.ZN(n2481));
   AOI22_X1 U3104 (.A1(REGISTERS[242]),
	.A2(FE_OFN113_n2768),
	.B1(REGISTERS[178]),
	.B2(FE_OFN11_n2767),
	.ZN(n2480));
   AND4_X1 U3105 (.A1(n2483),
	.A2(n2482),
	.A3(n2481),
	.A4(n2480),
	.ZN(n2495));
   AOI22_X1 U3106 (.A1(REGISTERS[850]),
	.A2(FE_OFN13_n2762),
	.B1(REGISTERS[786]),
	.B2(FE_OFN135_n2761),
	.ZN(n2487));
   AOI22_X1 U3107 (.A1(REGISTERS[978]),
	.A2(FE_OFN54_n2764),
	.B1(REGISTERS[914]),
	.B2(FE_OFN110_n2763),
	.ZN(n2486));
   AOI22_X1 U3108 (.A1(REGISTERS[882]),
	.A2(FE_OFN8_n2766),
	.B1(REGISTERS[818]),
	.B2(FE_OFN51_n2765),
	.ZN(n2485));
   AOI22_X1 U3109 (.A1(REGISTERS[1010]),
	.A2(FE_OFN113_n2768),
	.B1(REGISTERS[946]),
	.B2(FE_OFN11_n2767),
	.ZN(n2484));
   NAND4_X1 U3110 (.A1(n2487),
	.A2(n2486),
	.A3(n2485),
	.A4(n2484),
	.ZN(n2493));
   AOI22_X1 U3111 (.A1(REGISTERS[594]),
	.A2(FE_OFN13_n2762),
	.B1(REGISTERS[530]),
	.B2(FE_OFN135_n2761),
	.ZN(n2491));
   AOI22_X1 U3112 (.A1(REGISTERS[722]),
	.A2(FE_OFN54_n2764),
	.B1(REGISTERS[658]),
	.B2(FE_OFN110_n2763),
	.ZN(n2490));
   AOI22_X1 U3113 (.A1(REGISTERS[626]),
	.A2(FE_OFN8_n2766),
	.B1(REGISTERS[562]),
	.B2(FE_OFN51_n2765),
	.ZN(n2489));
   AOI22_X1 U3114 (.A1(REGISTERS[754]),
	.A2(FE_OFN113_n2768),
	.B1(REGISTERS[690]),
	.B2(FE_OFN11_n2767),
	.ZN(n2488));
   NAND4_X1 U3115 (.A1(n2491),
	.A2(n2490),
	.A3(n2489),
	.A4(n2488),
	.ZN(n2492));
   AOI22_X1 U3116 (.A1(n2493),
	.A2(FE_OFN32_n2776),
	.B1(n2492),
	.B2(FE_OFN30_n2774),
	.ZN(n2494));
   OAI221_X1 U3117 (.A(n2494),
	.B1(n2780),
	.B2(n2496),
	.C1(n2778),
	.C2(n2495),
	.ZN(N44));
   AOI22_X1 U3118 (.A1(REGISTERS[339]),
	.A2(FE_OFN14_n2762),
	.B1(REGISTERS[275]),
	.B2(FE_OFN136_n2761),
	.ZN(n2500));
   AOI22_X1 U3119 (.A1(REGISTERS[467]),
	.A2(FE_OFN55_n2764),
	.B1(REGISTERS[403]),
	.B2(FE_OFN111_n2763),
	.ZN(n2499));
   AOI22_X1 U3120 (.A1(REGISTERS[371]),
	.A2(FE_OFN9_n2766),
	.B1(REGISTERS[307]),
	.B2(FE_OFN52_n2765),
	.ZN(n2498));
   AOI22_X1 U3121 (.A1(REGISTERS[499]),
	.A2(FE_OFN114_n2768),
	.B1(REGISTERS[435]),
	.B2(FE_OFN11_n2767),
	.ZN(n2497));
   AND4_X1 U3122 (.A1(n2500),
	.A2(n2499),
	.A3(n2498),
	.A4(n2497),
	.ZN(n2517));
   AOI22_X1 U3123 (.A1(REGISTERS[83]),
	.A2(FE_OFN14_n2762),
	.B1(REGISTERS[19]),
	.B2(FE_OFN136_n2761),
	.ZN(n2504));
   AOI22_X1 U3124 (.A1(REGISTERS[211]),
	.A2(FE_OFN55_n2764),
	.B1(REGISTERS[147]),
	.B2(FE_OFN111_n2763),
	.ZN(n2503));
   AOI22_X1 U3125 (.A1(REGISTERS[115]),
	.A2(FE_OFN9_n2766),
	.B1(REGISTERS[51]),
	.B2(FE_OFN52_n2765),
	.ZN(n2502));
   AOI22_X1 U3126 (.A1(REGISTERS[243]),
	.A2(FE_OFN114_n2768),
	.B1(REGISTERS[179]),
	.B2(FE_OFN11_n2767),
	.ZN(n2501));
   AND4_X1 U3127 (.A1(n2504),
	.A2(n2503),
	.A3(n2502),
	.A4(n2501),
	.ZN(n2516));
   AOI22_X1 U3128 (.A1(REGISTERS[851]),
	.A2(FE_OFN14_n2762),
	.B1(REGISTERS[787]),
	.B2(FE_OFN136_n2761),
	.ZN(n2508));
   AOI22_X1 U3129 (.A1(REGISTERS[979]),
	.A2(FE_OFN56_n2764),
	.B1(REGISTERS[915]),
	.B2(FE_OFN112_n2763),
	.ZN(n2507));
   AOI22_X1 U3130 (.A1(REGISTERS[883]),
	.A2(FE_OFN10_n2766),
	.B1(REGISTERS[819]),
	.B2(FE_OFN53_n2765),
	.ZN(n2506));
   AOI22_X1 U3131 (.A1(REGISTERS[1011]),
	.A2(FE_OFN114_n2768),
	.B1(REGISTERS[947]),
	.B2(FE_OFN12_n2767),
	.ZN(n2505));
   NAND4_X1 U3132 (.A1(n2508),
	.A2(n2507),
	.A3(n2506),
	.A4(n2505),
	.ZN(n2514));
   AOI22_X1 U3133 (.A1(REGISTERS[595]),
	.A2(FE_OFN14_n2762),
	.B1(REGISTERS[531]),
	.B2(FE_OFN136_n2761),
	.ZN(n2512));
   AOI22_X1 U3134 (.A1(REGISTERS[723]),
	.A2(FE_OFN56_n2764),
	.B1(REGISTERS[659]),
	.B2(FE_OFN112_n2763),
	.ZN(n2511));
   AOI22_X1 U3135 (.A1(REGISTERS[627]),
	.A2(FE_OFN10_n2766),
	.B1(REGISTERS[563]),
	.B2(FE_OFN53_n2765),
	.ZN(n2510));
   AOI22_X1 U3136 (.A1(REGISTERS[755]),
	.A2(FE_OFN114_n2768),
	.B1(REGISTERS[691]),
	.B2(FE_OFN12_n2767),
	.ZN(n2509));
   NAND4_X1 U3137 (.A1(n2512),
	.A2(n2511),
	.A3(n2510),
	.A4(n2509),
	.ZN(n2513));
   AOI22_X1 U3138 (.A1(n2514),
	.A2(FE_OFN32_n2776),
	.B1(n2513),
	.B2(FE_OFN30_n2774),
	.ZN(n2515));
   OAI221_X1 U3139 (.A(n2515),
	.B1(n2780),
	.B2(n2517),
	.C1(n2778),
	.C2(n2516),
	.ZN(N43));
   AOI22_X1 U3140 (.A1(REGISTERS[340]),
	.A2(FE_OFN13_n2762),
	.B1(REGISTERS[276]),
	.B2(FE_OFN135_n2761),
	.ZN(n2521));
   AOI22_X1 U3141 (.A1(REGISTERS[468]),
	.A2(n2764),
	.B1(REGISTERS[404]),
	.B2(n2763),
	.ZN(n2520));
   AOI22_X1 U3142 (.A1(REGISTERS[372]),
	.A2(FE_OFN8_n2766),
	.B1(REGISTERS[308]),
	.B2(FE_OFN51_n2765),
	.ZN(n2519));
   AOI22_X1 U3143 (.A1(REGISTERS[500]),
	.A2(FE_OFN113_n2768),
	.B1(REGISTERS[436]),
	.B2(FE_OFN11_n2767),
	.ZN(n2518));
   AND4_X1 U3144 (.A1(n2521),
	.A2(n2520),
	.A3(n2519),
	.A4(n2518),
	.ZN(n2538));
   AOI22_X1 U3145 (.A1(REGISTERS[84]),
	.A2(FE_OFN13_n2762),
	.B1(REGISTERS[20]),
	.B2(FE_OFN135_n2761),
	.ZN(n2525));
   AOI22_X1 U3146 (.A1(REGISTERS[212]),
	.A2(n2764),
	.B1(REGISTERS[148]),
	.B2(n2763),
	.ZN(n2524));
   AOI22_X1 U3147 (.A1(REGISTERS[116]),
	.A2(FE_OFN8_n2766),
	.B1(REGISTERS[52]),
	.B2(FE_OFN51_n2765),
	.ZN(n2523));
   AOI22_X1 U3148 (.A1(REGISTERS[244]),
	.A2(FE_OFN113_n2768),
	.B1(REGISTERS[180]),
	.B2(FE_OFN11_n2767),
	.ZN(n2522));
   AND4_X1 U3149 (.A1(n2525),
	.A2(n2524),
	.A3(n2523),
	.A4(n2522),
	.ZN(n2537));
   AOI22_X1 U3150 (.A1(REGISTERS[852]),
	.A2(FE_OFN13_n2762),
	.B1(REGISTERS[788]),
	.B2(FE_OFN135_n2761),
	.ZN(n2529));
   AOI22_X1 U3151 (.A1(REGISTERS[980]),
	.A2(FE_OFN54_n2764),
	.B1(REGISTERS[916]),
	.B2(FE_OFN110_n2763),
	.ZN(n2528));
   AOI22_X1 U3152 (.A1(REGISTERS[884]),
	.A2(FE_OFN8_n2766),
	.B1(REGISTERS[820]),
	.B2(FE_OFN51_n2765),
	.ZN(n2527));
   AOI22_X1 U3153 (.A1(REGISTERS[1012]),
	.A2(FE_OFN113_n2768),
	.B1(REGISTERS[948]),
	.B2(FE_OFN11_n2767),
	.ZN(n2526));
   NAND4_X1 U3154 (.A1(n2529),
	.A2(n2528),
	.A3(n2527),
	.A4(n2526),
	.ZN(n2535));
   AOI22_X1 U3155 (.A1(REGISTERS[596]),
	.A2(FE_OFN13_n2762),
	.B1(REGISTERS[532]),
	.B2(FE_OFN135_n2761),
	.ZN(n2533));
   AOI22_X1 U3156 (.A1(REGISTERS[724]),
	.A2(FE_OFN54_n2764),
	.B1(REGISTERS[660]),
	.B2(FE_OFN110_n2763),
	.ZN(n2532));
   AOI22_X1 U3157 (.A1(REGISTERS[628]),
	.A2(FE_OFN8_n2766),
	.B1(REGISTERS[564]),
	.B2(FE_OFN51_n2765),
	.ZN(n2531));
   AOI22_X1 U3158 (.A1(REGISTERS[756]),
	.A2(FE_OFN113_n2768),
	.B1(REGISTERS[692]),
	.B2(FE_OFN11_n2767),
	.ZN(n2530));
   NAND4_X1 U3159 (.A1(n2533),
	.A2(n2532),
	.A3(n2531),
	.A4(n2530),
	.ZN(n2534));
   AOI22_X1 U3160 (.A1(n2535),
	.A2(FE_OFN32_n2776),
	.B1(n2534),
	.B2(FE_OFN30_n2774),
	.ZN(n2536));
   OAI221_X1 U3161 (.A(n2536),
	.B1(n2780),
	.B2(n2538),
	.C1(n2778),
	.C2(n2537),
	.ZN(N42));
   AOI22_X1 U3162 (.A1(REGISTERS[341]),
	.A2(FE_OFN13_n2762),
	.B1(REGISTERS[277]),
	.B2(FE_OFN135_n2761),
	.ZN(n2542));
   AOI22_X1 U3163 (.A1(REGISTERS[469]),
	.A2(FE_OFN55_n2764),
	.B1(REGISTERS[405]),
	.B2(FE_OFN112_n2763),
	.ZN(n2541));
   AOI22_X1 U3164 (.A1(REGISTERS[373]),
	.A2(FE_OFN8_n2766),
	.B1(REGISTERS[309]),
	.B2(FE_OFN51_n2765),
	.ZN(n2540));
   AOI22_X1 U3165 (.A1(REGISTERS[501]),
	.A2(FE_OFN113_n2768),
	.B1(REGISTERS[437]),
	.B2(FE_OFN11_n2767),
	.ZN(n2539));
   AND4_X1 U3166 (.A1(n2542),
	.A2(n2541),
	.A3(n2540),
	.A4(n2539),
	.ZN(n2559));
   AOI22_X1 U3167 (.A1(REGISTERS[85]),
	.A2(FE_OFN14_n2762),
	.B1(REGISTERS[21]),
	.B2(FE_OFN136_n2761),
	.ZN(n2546));
   AOI22_X1 U3168 (.A1(REGISTERS[213]),
	.A2(FE_OFN55_n2764),
	.B1(REGISTERS[149]),
	.B2(FE_OFN112_n2763),
	.ZN(n2545));
   AOI22_X1 U3169 (.A1(REGISTERS[117]),
	.A2(FE_OFN9_n2766),
	.B1(REGISTERS[53]),
	.B2(FE_OFN52_n2765),
	.ZN(n2544));
   AOI22_X1 U3170 (.A1(REGISTERS[245]),
	.A2(FE_OFN114_n2768),
	.B1(REGISTERS[181]),
	.B2(FE_OFN12_n2767),
	.ZN(n2543));
   AND4_X1 U3171 (.A1(n2546),
	.A2(n2545),
	.A3(n2544),
	.A4(n2543),
	.ZN(n2558));
   AOI22_X1 U3172 (.A1(REGISTERS[853]),
	.A2(FE_OFN14_n2762),
	.B1(REGISTERS[789]),
	.B2(FE_OFN136_n2761),
	.ZN(n2550));
   AOI22_X1 U3173 (.A1(REGISTERS[981]),
	.A2(FE_OFN55_n2764),
	.B1(REGISTERS[917]),
	.B2(FE_OFN112_n2763),
	.ZN(n2549));
   AOI22_X1 U3174 (.A1(REGISTERS[885]),
	.A2(FE_OFN9_n2766),
	.B1(REGISTERS[821]),
	.B2(FE_OFN52_n2765),
	.ZN(n2548));
   AOI22_X1 U3175 (.A1(REGISTERS[1013]),
	.A2(FE_OFN114_n2768),
	.B1(REGISTERS[949]),
	.B2(FE_OFN12_n2767),
	.ZN(n2547));
   NAND4_X1 U3176 (.A1(n2550),
	.A2(n2549),
	.A3(n2548),
	.A4(n2547),
	.ZN(n2556));
   AOI22_X1 U3177 (.A1(REGISTERS[597]),
	.A2(FE_OFN14_n2762),
	.B1(REGISTERS[533]),
	.B2(FE_OFN136_n2761),
	.ZN(n2554));
   AOI22_X1 U3178 (.A1(REGISTERS[725]),
	.A2(FE_OFN55_n2764),
	.B1(REGISTERS[661]),
	.B2(FE_OFN112_n2763),
	.ZN(n2553));
   AOI22_X1 U3179 (.A1(REGISTERS[629]),
	.A2(FE_OFN9_n2766),
	.B1(REGISTERS[565]),
	.B2(FE_OFN52_n2765),
	.ZN(n2552));
   AOI22_X1 U3180 (.A1(REGISTERS[757]),
	.A2(FE_OFN114_n2768),
	.B1(REGISTERS[693]),
	.B2(FE_OFN12_n2767),
	.ZN(n2551));
   NAND4_X1 U3181 (.A1(n2554),
	.A2(n2553),
	.A3(n2552),
	.A4(n2551),
	.ZN(n2555));
   AOI22_X1 U3182 (.A1(n2556),
	.A2(FE_OFN32_n2776),
	.B1(n2555),
	.B2(FE_OFN30_n2774),
	.ZN(n2557));
   OAI221_X1 U3183 (.A(n2557),
	.B1(n2780),
	.B2(n2559),
	.C1(n2778),
	.C2(n2558),
	.ZN(N41));
   AOI22_X1 U3184 (.A1(REGISTERS[342]),
	.A2(FE_OFN13_n2762),
	.B1(REGISTERS[278]),
	.B2(FE_OFN135_n2761),
	.ZN(n2563));
   AOI22_X1 U3185 (.A1(REGISTERS[470]),
	.A2(FE_OFN55_n2764),
	.B1(REGISTERS[406]),
	.B2(FE_OFN112_n2763),
	.ZN(n2562));
   AOI22_X1 U3186 (.A1(REGISTERS[374]),
	.A2(FE_OFN8_n2766),
	.B1(REGISTERS[310]),
	.B2(FE_OFN51_n2765),
	.ZN(n2561));
   AOI22_X1 U3187 (.A1(REGISTERS[502]),
	.A2(FE_OFN113_n2768),
	.B1(REGISTERS[438]),
	.B2(FE_OFN11_n2767),
	.ZN(n2560));
   AND4_X1 U3188 (.A1(n2563),
	.A2(n2562),
	.A3(n2561),
	.A4(n2560),
	.ZN(n2580));
   AOI22_X1 U3189 (.A1(REGISTERS[86]),
	.A2(FE_OFN13_n2762),
	.B1(REGISTERS[22]),
	.B2(FE_OFN135_n2761),
	.ZN(n2567));
   AOI22_X1 U3190 (.A1(REGISTERS[214]),
	.A2(FE_OFN55_n2764),
	.B1(REGISTERS[150]),
	.B2(FE_OFN112_n2763),
	.ZN(n2566));
   AOI22_X1 U3191 (.A1(REGISTERS[118]),
	.A2(FE_OFN8_n2766),
	.B1(REGISTERS[54]),
	.B2(FE_OFN51_n2765),
	.ZN(n2565));
   AOI22_X1 U3192 (.A1(REGISTERS[246]),
	.A2(FE_OFN113_n2768),
	.B1(REGISTERS[182]),
	.B2(FE_OFN11_n2767),
	.ZN(n2564));
   AND4_X1 U3193 (.A1(n2567),
	.A2(n2566),
	.A3(n2565),
	.A4(n2564),
	.ZN(n2579));
   AOI22_X1 U3194 (.A1(REGISTERS[854]),
	.A2(FE_OFN14_n2762),
	.B1(REGISTERS[790]),
	.B2(FE_OFN136_n2761),
	.ZN(n2571));
   AOI22_X1 U3195 (.A1(REGISTERS[982]),
	.A2(FE_OFN55_n2764),
	.B1(REGISTERS[918]),
	.B2(FE_OFN112_n2763),
	.ZN(n2570));
   AOI22_X1 U3196 (.A1(REGISTERS[886]),
	.A2(FE_OFN10_n2766),
	.B1(REGISTERS[822]),
	.B2(FE_OFN53_n2765),
	.ZN(n2569));
   AOI22_X1 U3197 (.A1(REGISTERS[1014]),
	.A2(FE_OFN114_n2768),
	.B1(REGISTERS[950]),
	.B2(FE_OFN12_n2767),
	.ZN(n2568));
   NAND4_X1 U3198 (.A1(n2571),
	.A2(n2570),
	.A3(n2569),
	.A4(n2568),
	.ZN(n2577));
   AOI22_X1 U3199 (.A1(REGISTERS[598]),
	.A2(FE_OFN14_n2762),
	.B1(REGISTERS[534]),
	.B2(FE_OFN136_n2761),
	.ZN(n2575));
   AOI22_X1 U3200 (.A1(REGISTERS[726]),
	.A2(FE_OFN55_n2764),
	.B1(REGISTERS[662]),
	.B2(FE_OFN112_n2763),
	.ZN(n2574));
   AOI22_X1 U3201 (.A1(REGISTERS[630]),
	.A2(FE_OFN10_n2766),
	.B1(REGISTERS[566]),
	.B2(FE_OFN53_n2765),
	.ZN(n2573));
   AOI22_X1 U3202 (.A1(REGISTERS[758]),
	.A2(FE_OFN114_n2768),
	.B1(REGISTERS[694]),
	.B2(FE_OFN12_n2767),
	.ZN(n2572));
   NAND4_X1 U3203 (.A1(n2575),
	.A2(n2574),
	.A3(n2573),
	.A4(n2572),
	.ZN(n2576));
   AOI22_X1 U3204 (.A1(n2577),
	.A2(FE_OFN32_n2776),
	.B1(n2576),
	.B2(FE_OFN30_n2774),
	.ZN(n2578));
   OAI221_X1 U3205 (.A(n2578),
	.B1(n2780),
	.B2(n2580),
	.C1(n2778),
	.C2(n2579),
	.ZN(N40));
   AOI22_X1 U3206 (.A1(REGISTERS[343]),
	.A2(FE_OFN14_n2762),
	.B1(REGISTERS[279]),
	.B2(FE_OFN136_n2761),
	.ZN(n2584));
   AOI22_X1 U3207 (.A1(REGISTERS[471]),
	.A2(FE_OFN55_n2764),
	.B1(REGISTERS[407]),
	.B2(FE_OFN111_n2763),
	.ZN(n2583));
   AOI22_X1 U3208 (.A1(REGISTERS[375]),
	.A2(FE_OFN9_n2766),
	.B1(REGISTERS[311]),
	.B2(FE_OFN52_n2765),
	.ZN(n2582));
   AOI22_X1 U3209 (.A1(REGISTERS[503]),
	.A2(FE_OFN114_n2768),
	.B1(REGISTERS[439]),
	.B2(FE_OFN11_n2767),
	.ZN(n2581));
   AND4_X1 U3210 (.A1(n2584),
	.A2(n2583),
	.A3(n2582),
	.A4(n2581),
	.ZN(n2601));
   AOI22_X1 U3211 (.A1(REGISTERS[87]),
	.A2(FE_OFN14_n2762),
	.B1(REGISTERS[23]),
	.B2(FE_OFN136_n2761),
	.ZN(n2588));
   AOI22_X1 U3212 (.A1(REGISTERS[215]),
	.A2(FE_OFN55_n2764),
	.B1(REGISTERS[151]),
	.B2(FE_OFN111_n2763),
	.ZN(n2587));
   AOI22_X1 U3213 (.A1(REGISTERS[119]),
	.A2(FE_OFN9_n2766),
	.B1(REGISTERS[55]),
	.B2(FE_OFN52_n2765),
	.ZN(n2586));
   AOI22_X1 U3214 (.A1(REGISTERS[247]),
	.A2(FE_OFN114_n2768),
	.B1(REGISTERS[183]),
	.B2(FE_OFN11_n2767),
	.ZN(n2585));
   AND4_X1 U3215 (.A1(n2588),
	.A2(n2587),
	.A3(n2586),
	.A4(n2585),
	.ZN(n2600));
   AOI22_X1 U3216 (.A1(REGISTERS[855]),
	.A2(FE_OFN14_n2762),
	.B1(REGISTERS[791]),
	.B2(FE_OFN136_n2761),
	.ZN(n2592));
   AOI22_X1 U3217 (.A1(REGISTERS[983]),
	.A2(FE_OFN55_n2764),
	.B1(REGISTERS[919]),
	.B2(FE_OFN112_n2763),
	.ZN(n2591));
   AOI22_X1 U3218 (.A1(REGISTERS[887]),
	.A2(FE_OFN10_n2766),
	.B1(REGISTERS[823]),
	.B2(FE_OFN53_n2765),
	.ZN(n2590));
   AOI22_X1 U3219 (.A1(REGISTERS[1015]),
	.A2(FE_OFN114_n2768),
	.B1(REGISTERS[951]),
	.B2(FE_OFN12_n2767),
	.ZN(n2589));
   NAND4_X1 U3220 (.A1(n2592),
	.A2(n2591),
	.A3(n2590),
	.A4(n2589),
	.ZN(n2598));
   AOI22_X1 U3221 (.A1(REGISTERS[599]),
	.A2(FE_OFN14_n2762),
	.B1(REGISTERS[535]),
	.B2(FE_OFN136_n2761),
	.ZN(n2596));
   AOI22_X1 U3222 (.A1(REGISTERS[727]),
	.A2(FE_OFN55_n2764),
	.B1(REGISTERS[663]),
	.B2(FE_OFN112_n2763),
	.ZN(n2595));
   AOI22_X1 U3223 (.A1(REGISTERS[631]),
	.A2(FE_OFN10_n2766),
	.B1(REGISTERS[567]),
	.B2(FE_OFN53_n2765),
	.ZN(n2594));
   AOI22_X1 U3224 (.A1(REGISTERS[759]),
	.A2(FE_OFN114_n2768),
	.B1(REGISTERS[695]),
	.B2(FE_OFN12_n2767),
	.ZN(n2593));
   NAND4_X1 U3225 (.A1(n2596),
	.A2(n2595),
	.A3(n2594),
	.A4(n2593),
	.ZN(n2597));
   AOI22_X1 U3226 (.A1(n2598),
	.A2(FE_OFN32_n2776),
	.B1(n2597),
	.B2(FE_OFN30_n2774),
	.ZN(n2599));
   OAI221_X1 U3227 (.A(n2599),
	.B1(n2780),
	.B2(n2601),
	.C1(n2778),
	.C2(n2600),
	.ZN(N39));
   AOI22_X1 U3228 (.A1(REGISTERS[344]),
	.A2(FE_OFN13_n2762),
	.B1(REGISTERS[280]),
	.B2(FE_OFN135_n2761),
	.ZN(n2605));
   AOI22_X1 U3229 (.A1(REGISTERS[472]),
	.A2(n2764),
	.B1(REGISTERS[408]),
	.B2(n2763),
	.ZN(n2604));
   AOI22_X1 U3230 (.A1(REGISTERS[376]),
	.A2(FE_OFN8_n2766),
	.B1(REGISTERS[312]),
	.B2(FE_OFN51_n2765),
	.ZN(n2603));
   AOI22_X1 U3231 (.A1(REGISTERS[504]),
	.A2(FE_OFN113_n2768),
	.B1(REGISTERS[440]),
	.B2(FE_OFN11_n2767),
	.ZN(n2602));
   AND4_X1 U3232 (.A1(n2605),
	.A2(n2604),
	.A3(n2603),
	.A4(n2602),
	.ZN(n2622));
   AOI22_X1 U3233 (.A1(REGISTERS[88]),
	.A2(FE_OFN13_n2762),
	.B1(REGISTERS[24]),
	.B2(FE_OFN135_n2761),
	.ZN(n2609));
   AOI22_X1 U3234 (.A1(REGISTERS[216]),
	.A2(n2764),
	.B1(REGISTERS[152]),
	.B2(n2763),
	.ZN(n2608));
   AOI22_X1 U3235 (.A1(REGISTERS[120]),
	.A2(FE_OFN8_n2766),
	.B1(REGISTERS[56]),
	.B2(FE_OFN51_n2765),
	.ZN(n2607));
   AOI22_X1 U3236 (.A1(REGISTERS[248]),
	.A2(FE_OFN113_n2768),
	.B1(REGISTERS[184]),
	.B2(FE_OFN11_n2767),
	.ZN(n2606));
   AND4_X1 U3237 (.A1(n2609),
	.A2(n2608),
	.A3(n2607),
	.A4(n2606),
	.ZN(n2621));
   AOI22_X1 U3238 (.A1(REGISTERS[856]),
	.A2(FE_OFN13_n2762),
	.B1(REGISTERS[792]),
	.B2(FE_OFN135_n2761),
	.ZN(n2613));
   AOI22_X1 U3239 (.A1(REGISTERS[984]),
	.A2(FE_OFN54_n2764),
	.B1(REGISTERS[920]),
	.B2(FE_OFN110_n2763),
	.ZN(n2612));
   AOI22_X1 U3240 (.A1(REGISTERS[888]),
	.A2(FE_OFN8_n2766),
	.B1(REGISTERS[824]),
	.B2(FE_OFN51_n2765),
	.ZN(n2611));
   AOI22_X1 U3241 (.A1(REGISTERS[1016]),
	.A2(FE_OFN113_n2768),
	.B1(REGISTERS[952]),
	.B2(FE_OFN11_n2767),
	.ZN(n2610));
   NAND4_X1 U3242 (.A1(n2613),
	.A2(n2612),
	.A3(n2611),
	.A4(n2610),
	.ZN(n2619));
   AOI22_X1 U3243 (.A1(REGISTERS[600]),
	.A2(FE_OFN13_n2762),
	.B1(REGISTERS[536]),
	.B2(FE_OFN135_n2761),
	.ZN(n2617));
   AOI22_X1 U3244 (.A1(REGISTERS[728]),
	.A2(FE_OFN54_n2764),
	.B1(REGISTERS[664]),
	.B2(FE_OFN110_n2763),
	.ZN(n2616));
   AOI22_X1 U3245 (.A1(REGISTERS[632]),
	.A2(FE_OFN8_n2766),
	.B1(REGISTERS[568]),
	.B2(FE_OFN51_n2765),
	.ZN(n2615));
   AOI22_X1 U3246 (.A1(REGISTERS[760]),
	.A2(FE_OFN113_n2768),
	.B1(REGISTERS[696]),
	.B2(FE_OFN11_n2767),
	.ZN(n2614));
   NAND4_X1 U3247 (.A1(n2617),
	.A2(n2616),
	.A3(n2615),
	.A4(n2614),
	.ZN(n2618));
   AOI22_X1 U3248 (.A1(n2619),
	.A2(FE_OFN32_n2776),
	.B1(n2618),
	.B2(FE_OFN30_n2774),
	.ZN(n2620));
   OAI221_X1 U3249 (.A(n2620),
	.B1(n2780),
	.B2(n2622),
	.C1(n2778),
	.C2(n2621),
	.ZN(N38));
   AOI22_X1 U3250 (.A1(REGISTERS[345]),
	.A2(FE_OFN14_n2762),
	.B1(REGISTERS[281]),
	.B2(FE_OFN136_n2761),
	.ZN(n2626));
   AOI22_X1 U3251 (.A1(REGISTERS[473]),
	.A2(FE_OFN55_n2764),
	.B1(REGISTERS[409]),
	.B2(FE_OFN111_n2763),
	.ZN(n2625));
   AOI22_X1 U3252 (.A1(REGISTERS[377]),
	.A2(FE_OFN9_n2766),
	.B1(REGISTERS[313]),
	.B2(FE_OFN52_n2765),
	.ZN(n2624));
   AOI22_X1 U3253 (.A1(REGISTERS[505]),
	.A2(FE_OFN114_n2768),
	.B1(REGISTERS[441]),
	.B2(FE_OFN11_n2767),
	.ZN(n2623));
   AND4_X1 U3254 (.A1(n2626),
	.A2(n2625),
	.A3(n2624),
	.A4(n2623),
	.ZN(n2643));
   AOI22_X1 U3255 (.A1(REGISTERS[89]),
	.A2(FE_OFN14_n2762),
	.B1(REGISTERS[25]),
	.B2(FE_OFN136_n2761),
	.ZN(n2630));
   AOI22_X1 U3256 (.A1(REGISTERS[217]),
	.A2(FE_OFN55_n2764),
	.B1(REGISTERS[153]),
	.B2(FE_OFN111_n2763),
	.ZN(n2629));
   AOI22_X1 U3257 (.A1(REGISTERS[121]),
	.A2(FE_OFN9_n2766),
	.B1(REGISTERS[57]),
	.B2(FE_OFN52_n2765),
	.ZN(n2628));
   AOI22_X1 U3258 (.A1(REGISTERS[249]),
	.A2(FE_OFN114_n2768),
	.B1(REGISTERS[185]),
	.B2(FE_OFN11_n2767),
	.ZN(n2627));
   AND4_X1 U3259 (.A1(n2630),
	.A2(n2629),
	.A3(n2628),
	.A4(n2627),
	.ZN(n2642));
   AOI22_X1 U3260 (.A1(REGISTERS[857]),
	.A2(FE_OFN14_n2762),
	.B1(REGISTERS[793]),
	.B2(FE_OFN136_n2761),
	.ZN(n2634));
   AOI22_X1 U3261 (.A1(REGISTERS[985]),
	.A2(FE_OFN55_n2764),
	.B1(REGISTERS[921]),
	.B2(FE_OFN112_n2763),
	.ZN(n2633));
   AOI22_X1 U3262 (.A1(REGISTERS[889]),
	.A2(FE_OFN10_n2766),
	.B1(REGISTERS[825]),
	.B2(FE_OFN53_n2765),
	.ZN(n2632));
   AOI22_X1 U3263 (.A1(REGISTERS[1017]),
	.A2(FE_OFN114_n2768),
	.B1(REGISTERS[953]),
	.B2(FE_OFN12_n2767),
	.ZN(n2631));
   NAND4_X1 U3264 (.A1(n2634),
	.A2(n2633),
	.A3(n2632),
	.A4(n2631),
	.ZN(n2640));
   AOI22_X1 U3265 (.A1(REGISTERS[601]),
	.A2(FE_OFN14_n2762),
	.B1(REGISTERS[537]),
	.B2(FE_OFN136_n2761),
	.ZN(n2638));
   AOI22_X1 U3266 (.A1(REGISTERS[729]),
	.A2(FE_OFN55_n2764),
	.B1(REGISTERS[665]),
	.B2(FE_OFN112_n2763),
	.ZN(n2637));
   AOI22_X1 U3267 (.A1(REGISTERS[633]),
	.A2(FE_OFN10_n2766),
	.B1(REGISTERS[569]),
	.B2(FE_OFN53_n2765),
	.ZN(n2636));
   AOI22_X1 U3268 (.A1(REGISTERS[761]),
	.A2(FE_OFN114_n2768),
	.B1(REGISTERS[697]),
	.B2(FE_OFN12_n2767),
	.ZN(n2635));
   NAND4_X1 U3269 (.A1(n2638),
	.A2(n2637),
	.A3(n2636),
	.A4(n2635),
	.ZN(n2639));
   AOI22_X1 U3270 (.A1(n2640),
	.A2(FE_OFN32_n2776),
	.B1(n2639),
	.B2(FE_OFN30_n2774),
	.ZN(n2641));
   OAI221_X1 U3271 (.A(n2641),
	.B1(n2780),
	.B2(n2643),
	.C1(n2778),
	.C2(n2642),
	.ZN(N37));
   AOI22_X1 U3272 (.A1(REGISTERS[346]),
	.A2(FE_OFN13_n2762),
	.B1(REGISTERS[282]),
	.B2(FE_OFN135_n2761),
	.ZN(n2647));
   AOI22_X1 U3273 (.A1(REGISTERS[474]),
	.A2(n2764),
	.B1(REGISTERS[410]),
	.B2(n2763),
	.ZN(n2646));
   AOI22_X1 U3274 (.A1(REGISTERS[378]),
	.A2(FE_OFN8_n2766),
	.B1(REGISTERS[314]),
	.B2(FE_OFN51_n2765),
	.ZN(n2645));
   AOI22_X1 U3275 (.A1(REGISTERS[506]),
	.A2(FE_OFN113_n2768),
	.B1(REGISTERS[442]),
	.B2(FE_OFN11_n2767),
	.ZN(n2644));
   AND4_X1 U3276 (.A1(n2647),
	.A2(n2646),
	.A3(n2645),
	.A4(n2644),
	.ZN(n2664));
   AOI22_X1 U3277 (.A1(REGISTERS[90]),
	.A2(FE_OFN13_n2762),
	.B1(REGISTERS[26]),
	.B2(FE_OFN135_n2761),
	.ZN(n2651));
   AOI22_X1 U3278 (.A1(REGISTERS[218]),
	.A2(n2764),
	.B1(REGISTERS[154]),
	.B2(n2763),
	.ZN(n2650));
   AOI22_X1 U3279 (.A1(REGISTERS[122]),
	.A2(FE_OFN8_n2766),
	.B1(REGISTERS[58]),
	.B2(FE_OFN51_n2765),
	.ZN(n2649));
   AOI22_X1 U3280 (.A1(REGISTERS[250]),
	.A2(FE_OFN113_n2768),
	.B1(REGISTERS[186]),
	.B2(FE_OFN11_n2767),
	.ZN(n2648));
   AND4_X1 U3281 (.A1(n2651),
	.A2(n2650),
	.A3(n2649),
	.A4(n2648),
	.ZN(n2663));
   AOI22_X1 U3282 (.A1(REGISTERS[858]),
	.A2(FE_OFN13_n2762),
	.B1(REGISTERS[794]),
	.B2(FE_OFN135_n2761),
	.ZN(n2655));
   AOI22_X1 U3283 (.A1(REGISTERS[986]),
	.A2(FE_OFN54_n2764),
	.B1(REGISTERS[922]),
	.B2(FE_OFN110_n2763),
	.ZN(n2654));
   AOI22_X1 U3284 (.A1(REGISTERS[890]),
	.A2(FE_OFN8_n2766),
	.B1(REGISTERS[826]),
	.B2(FE_OFN51_n2765),
	.ZN(n2653));
   AOI22_X1 U3285 (.A1(REGISTERS[1018]),
	.A2(FE_OFN113_n2768),
	.B1(REGISTERS[954]),
	.B2(FE_OFN11_n2767),
	.ZN(n2652));
   NAND4_X1 U3286 (.A1(n2655),
	.A2(n2654),
	.A3(n2653),
	.A4(n2652),
	.ZN(n2661));
   AOI22_X1 U3287 (.A1(REGISTERS[602]),
	.A2(FE_OFN13_n2762),
	.B1(REGISTERS[538]),
	.B2(FE_OFN135_n2761),
	.ZN(n2659));
   AOI22_X1 U3288 (.A1(REGISTERS[730]),
	.A2(FE_OFN54_n2764),
	.B1(REGISTERS[666]),
	.B2(FE_OFN110_n2763),
	.ZN(n2658));
   AOI22_X1 U3289 (.A1(REGISTERS[634]),
	.A2(FE_OFN8_n2766),
	.B1(REGISTERS[570]),
	.B2(FE_OFN51_n2765),
	.ZN(n2657));
   AOI22_X1 U3290 (.A1(REGISTERS[762]),
	.A2(FE_OFN113_n2768),
	.B1(REGISTERS[698]),
	.B2(FE_OFN11_n2767),
	.ZN(n2656));
   NAND4_X1 U3291 (.A1(n2659),
	.A2(n2658),
	.A3(n2657),
	.A4(n2656),
	.ZN(n2660));
   AOI22_X1 U3292 (.A1(n2661),
	.A2(FE_OFN32_n2776),
	.B1(n2660),
	.B2(FE_OFN30_n2774),
	.ZN(n2662));
   OAI221_X1 U3293 (.A(n2662),
	.B1(n2780),
	.B2(n2664),
	.C1(n2778),
	.C2(n2663),
	.ZN(N36));
   AOI22_X1 U3294 (.A1(REGISTERS[347]),
	.A2(FE_OFN14_n2762),
	.B1(REGISTERS[283]),
	.B2(FE_OFN136_n2761),
	.ZN(n2668));
   AOI22_X1 U3295 (.A1(REGISTERS[475]),
	.A2(FE_OFN55_n2764),
	.B1(REGISTERS[411]),
	.B2(FE_OFN111_n2763),
	.ZN(n2667));
   AOI22_X1 U3296 (.A1(REGISTERS[379]),
	.A2(FE_OFN9_n2766),
	.B1(REGISTERS[315]),
	.B2(FE_OFN52_n2765),
	.ZN(n2666));
   AOI22_X1 U3297 (.A1(REGISTERS[507]),
	.A2(FE_OFN114_n2768),
	.B1(REGISTERS[443]),
	.B2(FE_OFN12_n2767),
	.ZN(n2665));
   AND4_X1 U3298 (.A1(n2668),
	.A2(n2667),
	.A3(n2666),
	.A4(n2665),
	.ZN(n2685));
   AOI22_X1 U3299 (.A1(REGISTERS[91]),
	.A2(FE_OFN14_n2762),
	.B1(REGISTERS[27]),
	.B2(FE_OFN136_n2761),
	.ZN(n2672));
   AOI22_X1 U3300 (.A1(REGISTERS[219]),
	.A2(FE_OFN55_n2764),
	.B1(REGISTERS[155]),
	.B2(FE_OFN111_n2763),
	.ZN(n2671));
   AOI22_X1 U3301 (.A1(REGISTERS[123]),
	.A2(FE_OFN9_n2766),
	.B1(REGISTERS[59]),
	.B2(FE_OFN52_n2765),
	.ZN(n2670));
   AOI22_X1 U3302 (.A1(REGISTERS[251]),
	.A2(FE_OFN114_n2768),
	.B1(REGISTERS[187]),
	.B2(FE_OFN12_n2767),
	.ZN(n2669));
   AND4_X1 U3303 (.A1(n2672),
	.A2(n2671),
	.A3(n2670),
	.A4(n2669),
	.ZN(n2684));
   AOI22_X1 U3304 (.A1(REGISTERS[859]),
	.A2(FE_OFN14_n2762),
	.B1(REGISTERS[795]),
	.B2(FE_OFN136_n2761),
	.ZN(n2676));
   AOI22_X1 U3305 (.A1(REGISTERS[987]),
	.A2(FE_OFN56_n2764),
	.B1(REGISTERS[923]),
	.B2(FE_OFN112_n2763),
	.ZN(n2675));
   AOI22_X1 U3306 (.A1(REGISTERS[891]),
	.A2(FE_OFN10_n2766),
	.B1(REGISTERS[827]),
	.B2(FE_OFN53_n2765),
	.ZN(n2674));
   AOI22_X1 U3307 (.A1(REGISTERS[1019]),
	.A2(FE_OFN114_n2768),
	.B1(REGISTERS[955]),
	.B2(FE_OFN12_n2767),
	.ZN(n2673));
   NAND4_X1 U3308 (.A1(n2676),
	.A2(n2675),
	.A3(n2674),
	.A4(n2673),
	.ZN(n2682));
   AOI22_X1 U3309 (.A1(REGISTERS[603]),
	.A2(FE_OFN14_n2762),
	.B1(REGISTERS[539]),
	.B2(FE_OFN136_n2761),
	.ZN(n2680));
   AOI22_X1 U3310 (.A1(REGISTERS[731]),
	.A2(FE_OFN56_n2764),
	.B1(REGISTERS[667]),
	.B2(FE_OFN112_n2763),
	.ZN(n2679));
   AOI22_X1 U3311 (.A1(REGISTERS[635]),
	.A2(FE_OFN10_n2766),
	.B1(REGISTERS[571]),
	.B2(FE_OFN53_n2765),
	.ZN(n2678));
   AOI22_X1 U3312 (.A1(REGISTERS[763]),
	.A2(FE_OFN114_n2768),
	.B1(REGISTERS[699]),
	.B2(FE_OFN12_n2767),
	.ZN(n2677));
   NAND4_X1 U3313 (.A1(n2680),
	.A2(n2679),
	.A3(n2678),
	.A4(n2677),
	.ZN(n2681));
   AOI22_X1 U3314 (.A1(n2682),
	.A2(FE_OFN32_n2776),
	.B1(n2681),
	.B2(FE_OFN30_n2774),
	.ZN(n2683));
   OAI221_X1 U3315 (.A(n2683),
	.B1(n2780),
	.B2(n2685),
	.C1(n2778),
	.C2(n2684),
	.ZN(N35));
   AOI22_X1 U3316 (.A1(REGISTERS[348]),
	.A2(FE_OFN13_n2762),
	.B1(REGISTERS[284]),
	.B2(FE_OFN135_n2761),
	.ZN(n2689));
   AOI22_X1 U3317 (.A1(REGISTERS[476]),
	.A2(FE_OFN55_n2764),
	.B1(REGISTERS[412]),
	.B2(FE_OFN112_n2763),
	.ZN(n2688));
   AOI22_X1 U3318 (.A1(REGISTERS[380]),
	.A2(FE_OFN8_n2766),
	.B1(REGISTERS[316]),
	.B2(FE_OFN51_n2765),
	.ZN(n2687));
   AOI22_X1 U3319 (.A1(REGISTERS[508]),
	.A2(FE_OFN113_n2768),
	.B1(REGISTERS[444]),
	.B2(FE_OFN11_n2767),
	.ZN(n2686));
   AND4_X1 U3320 (.A1(n2689),
	.A2(n2688),
	.A3(n2687),
	.A4(n2686),
	.ZN(n2706));
   AOI22_X1 U3321 (.A1(REGISTERS[92]),
	.A2(FE_OFN13_n2762),
	.B1(REGISTERS[28]),
	.B2(FE_OFN135_n2761),
	.ZN(n2693));
   AOI22_X1 U3322 (.A1(REGISTERS[220]),
	.A2(FE_OFN55_n2764),
	.B1(REGISTERS[156]),
	.B2(FE_OFN112_n2763),
	.ZN(n2692));
   AOI22_X1 U3323 (.A1(REGISTERS[124]),
	.A2(FE_OFN8_n2766),
	.B1(REGISTERS[60]),
	.B2(FE_OFN51_n2765),
	.ZN(n2691));
   AOI22_X1 U3324 (.A1(REGISTERS[252]),
	.A2(FE_OFN113_n2768),
	.B1(REGISTERS[188]),
	.B2(FE_OFN11_n2767),
	.ZN(n2690));
   AND4_X1 U3325 (.A1(n2693),
	.A2(n2692),
	.A3(n2691),
	.A4(n2690),
	.ZN(n2705));
   AOI22_X1 U3326 (.A1(REGISTERS[860]),
	.A2(FE_OFN14_n2762),
	.B1(REGISTERS[796]),
	.B2(FE_OFN136_n2761),
	.ZN(n2697));
   AOI22_X1 U3327 (.A1(REGISTERS[988]),
	.A2(FE_OFN55_n2764),
	.B1(REGISTERS[924]),
	.B2(FE_OFN112_n2763),
	.ZN(n2696));
   AOI22_X1 U3328 (.A1(REGISTERS[892]),
	.A2(FE_OFN10_n2766),
	.B1(REGISTERS[828]),
	.B2(FE_OFN53_n2765),
	.ZN(n2695));
   AOI22_X1 U3329 (.A1(REGISTERS[1020]),
	.A2(FE_OFN114_n2768),
	.B1(REGISTERS[956]),
	.B2(FE_OFN12_n2767),
	.ZN(n2694));
   NAND4_X1 U3330 (.A1(n2697),
	.A2(n2696),
	.A3(n2695),
	.A4(n2694),
	.ZN(n2703));
   AOI22_X1 U3331 (.A1(REGISTERS[604]),
	.A2(FE_OFN14_n2762),
	.B1(REGISTERS[540]),
	.B2(FE_OFN136_n2761),
	.ZN(n2701));
   AOI22_X1 U3332 (.A1(REGISTERS[732]),
	.A2(FE_OFN55_n2764),
	.B1(REGISTERS[668]),
	.B2(FE_OFN112_n2763),
	.ZN(n2700));
   AOI22_X1 U3333 (.A1(REGISTERS[636]),
	.A2(FE_OFN10_n2766),
	.B1(REGISTERS[572]),
	.B2(FE_OFN53_n2765),
	.ZN(n2699));
   AOI22_X1 U3334 (.A1(REGISTERS[764]),
	.A2(FE_OFN114_n2768),
	.B1(REGISTERS[700]),
	.B2(FE_OFN12_n2767),
	.ZN(n2698));
   NAND4_X1 U3335 (.A1(n2701),
	.A2(n2700),
	.A3(n2699),
	.A4(n2698),
	.ZN(n2702));
   AOI22_X1 U3336 (.A1(n2703),
	.A2(FE_OFN32_n2776),
	.B1(n2702),
	.B2(FE_OFN30_n2774),
	.ZN(n2704));
   OAI221_X1 U3337 (.A(n2704),
	.B1(n2780),
	.B2(n2706),
	.C1(n2778),
	.C2(n2705),
	.ZN(N34));
   AOI22_X1 U3338 (.A1(REGISTERS[349]),
	.A2(FE_OFN13_n2762),
	.B1(REGISTERS[285]),
	.B2(FE_OFN135_n2761),
	.ZN(n2710));
   AOI22_X1 U3339 (.A1(REGISTERS[477]),
	.A2(FE_OFN54_n2764),
	.B1(REGISTERS[413]),
	.B2(FE_OFN110_n2763),
	.ZN(n2709));
   AOI22_X1 U3340 (.A1(REGISTERS[381]),
	.A2(FE_OFN8_n2766),
	.B1(REGISTERS[317]),
	.B2(n2765),
	.ZN(n2708));
   AOI22_X1 U3341 (.A1(REGISTERS[509]),
	.A2(FE_OFN113_n2768),
	.B1(REGISTERS[445]),
	.B2(FE_OFN11_n2767),
	.ZN(n2707));
   AND4_X1 U3342 (.A1(n2710),
	.A2(n2709),
	.A3(n2708),
	.A4(n2707),
	.ZN(n2727));
   AOI22_X1 U3343 (.A1(REGISTERS[93]),
	.A2(FE_OFN13_n2762),
	.B1(REGISTERS[29]),
	.B2(FE_OFN135_n2761),
	.ZN(n2714));
   AOI22_X1 U3344 (.A1(REGISTERS[221]),
	.A2(FE_OFN54_n2764),
	.B1(REGISTERS[157]),
	.B2(FE_OFN110_n2763),
	.ZN(n2713));
   AOI22_X1 U3345 (.A1(REGISTERS[125]),
	.A2(FE_OFN8_n2766),
	.B1(REGISTERS[61]),
	.B2(n2765),
	.ZN(n2712));
   AOI22_X1 U3346 (.A1(REGISTERS[253]),
	.A2(FE_OFN113_n2768),
	.B1(REGISTERS[189]),
	.B2(FE_OFN11_n2767),
	.ZN(n2711));
   AND4_X1 U3347 (.A1(n2714),
	.A2(n2713),
	.A3(n2712),
	.A4(n2711),
	.ZN(n2726));
   AOI22_X1 U3348 (.A1(REGISTERS[861]),
	.A2(FE_OFN13_n2762),
	.B1(REGISTERS[797]),
	.B2(FE_OFN135_n2761),
	.ZN(n2718));
   AOI22_X1 U3349 (.A1(REGISTERS[989]),
	.A2(FE_OFN54_n2764),
	.B1(REGISTERS[925]),
	.B2(FE_OFN110_n2763),
	.ZN(n2717));
   AOI22_X1 U3350 (.A1(REGISTERS[893]),
	.A2(FE_OFN8_n2766),
	.B1(REGISTERS[829]),
	.B2(FE_OFN51_n2765),
	.ZN(n2716));
   AOI22_X1 U3351 (.A1(REGISTERS[1021]),
	.A2(FE_OFN113_n2768),
	.B1(REGISTERS[957]),
	.B2(FE_OFN11_n2767),
	.ZN(n2715));
   NAND4_X1 U3352 (.A1(n2718),
	.A2(n2717),
	.A3(n2716),
	.A4(n2715),
	.ZN(n2724));
   AOI22_X1 U3353 (.A1(REGISTERS[605]),
	.A2(FE_OFN13_n2762),
	.B1(REGISTERS[541]),
	.B2(FE_OFN135_n2761),
	.ZN(n2722));
   AOI22_X1 U3354 (.A1(REGISTERS[733]),
	.A2(FE_OFN54_n2764),
	.B1(REGISTERS[669]),
	.B2(FE_OFN110_n2763),
	.ZN(n2721));
   AOI22_X1 U3355 (.A1(REGISTERS[637]),
	.A2(FE_OFN8_n2766),
	.B1(REGISTERS[573]),
	.B2(FE_OFN51_n2765),
	.ZN(n2720));
   AOI22_X1 U3356 (.A1(REGISTERS[765]),
	.A2(FE_OFN113_n2768),
	.B1(REGISTERS[701]),
	.B2(FE_OFN11_n2767),
	.ZN(n2719));
   NAND4_X1 U3357 (.A1(n2722),
	.A2(n2721),
	.A3(n2720),
	.A4(n2719),
	.ZN(n2723));
   AOI22_X1 U3358 (.A1(n2724),
	.A2(FE_OFN32_n2776),
	.B1(n2723),
	.B2(FE_OFN30_n2774),
	.ZN(n2725));
   OAI221_X1 U3359 (.A(n2725),
	.B1(n2780),
	.B2(n2727),
	.C1(n2778),
	.C2(n2726),
	.ZN(N33));
   AOI22_X1 U3360 (.A1(REGISTERS[350]),
	.A2(FE_OFN13_n2762),
	.B1(REGISTERS[286]),
	.B2(FE_OFN135_n2761),
	.ZN(n2731));
   AOI22_X1 U3361 (.A1(REGISTERS[478]),
	.A2(FE_OFN55_n2764),
	.B1(REGISTERS[414]),
	.B2(FE_OFN112_n2763),
	.ZN(n2730));
   AOI22_X1 U3362 (.A1(REGISTERS[382]),
	.A2(FE_OFN8_n2766),
	.B1(REGISTERS[318]),
	.B2(FE_OFN51_n2765),
	.ZN(n2729));
   AOI22_X1 U3363 (.A1(REGISTERS[510]),
	.A2(FE_OFN113_n2768),
	.B1(REGISTERS[446]),
	.B2(FE_OFN11_n2767),
	.ZN(n2728));
   AND4_X1 U3364 (.A1(n2731),
	.A2(n2730),
	.A3(n2729),
	.A4(n2728),
	.ZN(n2748));
   AOI22_X1 U3365 (.A1(REGISTERS[94]),
	.A2(FE_OFN13_n2762),
	.B1(REGISTERS[30]),
	.B2(FE_OFN135_n2761),
	.ZN(n2735));
   AOI22_X1 U3366 (.A1(REGISTERS[222]),
	.A2(FE_OFN55_n2764),
	.B1(REGISTERS[158]),
	.B2(FE_OFN112_n2763),
	.ZN(n2734));
   AOI22_X1 U3367 (.A1(REGISTERS[126]),
	.A2(FE_OFN8_n2766),
	.B1(REGISTERS[62]),
	.B2(FE_OFN51_n2765),
	.ZN(n2733));
   AOI22_X1 U3368 (.A1(REGISTERS[254]),
	.A2(FE_OFN113_n2768),
	.B1(REGISTERS[190]),
	.B2(FE_OFN11_n2767),
	.ZN(n2732));
   AND4_X1 U3369 (.A1(n2735),
	.A2(n2734),
	.A3(n2733),
	.A4(n2732),
	.ZN(n2747));
   AOI22_X1 U3370 (.A1(REGISTERS[862]),
	.A2(FE_OFN14_n2762),
	.B1(REGISTERS[798]),
	.B2(FE_OFN136_n2761),
	.ZN(n2739));
   AOI22_X1 U3371 (.A1(REGISTERS[990]),
	.A2(FE_OFN55_n2764),
	.B1(REGISTERS[926]),
	.B2(FE_OFN112_n2763),
	.ZN(n2738));
   AOI22_X1 U3372 (.A1(REGISTERS[894]),
	.A2(FE_OFN9_n2766),
	.B1(REGISTERS[830]),
	.B2(FE_OFN52_n2765),
	.ZN(n2737));
   AOI22_X1 U3373 (.A1(REGISTERS[1022]),
	.A2(FE_OFN114_n2768),
	.B1(REGISTERS[958]),
	.B2(FE_OFN12_n2767),
	.ZN(n2736));
   NAND4_X1 U3374 (.A1(n2739),
	.A2(n2738),
	.A3(n2737),
	.A4(n2736),
	.ZN(n2745));
   AOI22_X1 U3375 (.A1(REGISTERS[606]),
	.A2(FE_OFN14_n2762),
	.B1(REGISTERS[542]),
	.B2(FE_OFN136_n2761),
	.ZN(n2743));
   AOI22_X1 U3376 (.A1(REGISTERS[734]),
	.A2(FE_OFN55_n2764),
	.B1(REGISTERS[670]),
	.B2(FE_OFN112_n2763),
	.ZN(n2742));
   AOI22_X1 U3377 (.A1(REGISTERS[638]),
	.A2(FE_OFN9_n2766),
	.B1(REGISTERS[574]),
	.B2(FE_OFN52_n2765),
	.ZN(n2741));
   AOI22_X1 U3378 (.A1(REGISTERS[766]),
	.A2(FE_OFN114_n2768),
	.B1(REGISTERS[702]),
	.B2(FE_OFN12_n2767),
	.ZN(n2740));
   NAND4_X1 U3379 (.A1(n2743),
	.A2(n2742),
	.A3(n2741),
	.A4(n2740),
	.ZN(n2744));
   AOI22_X1 U3380 (.A1(n2745),
	.A2(FE_OFN32_n2776),
	.B1(n2744),
	.B2(FE_OFN30_n2774),
	.ZN(n2746));
   OAI221_X1 U3381 (.A(n2746),
	.B1(n2780),
	.B2(n2748),
	.C1(n2778),
	.C2(n2747),
	.ZN(N32));
   AOI22_X1 U3382 (.A1(REGISTERS[351]),
	.A2(FE_OFN13_n2762),
	.B1(REGISTERS[287]),
	.B2(FE_OFN135_n2761),
	.ZN(n2752));
   AOI22_X1 U3383 (.A1(REGISTERS[479]),
	.A2(n2764),
	.B1(REGISTERS[415]),
	.B2(n2763),
	.ZN(n2751));
   AOI22_X1 U3384 (.A1(REGISTERS[383]),
	.A2(FE_OFN8_n2766),
	.B1(REGISTERS[319]),
	.B2(FE_OFN51_n2765),
	.ZN(n2750));
   AOI22_X1 U3385 (.A1(REGISTERS[511]),
	.A2(FE_OFN113_n2768),
	.B1(REGISTERS[447]),
	.B2(FE_OFN11_n2767),
	.ZN(n2749));
   AND4_X1 U3386 (.A1(n2752),
	.A2(n2751),
	.A3(n2750),
	.A4(n2749),
	.ZN(n2781));
   AOI22_X1 U3387 (.A1(REGISTERS[95]),
	.A2(FE_OFN13_n2762),
	.B1(REGISTERS[31]),
	.B2(FE_OFN135_n2761),
	.ZN(n2756));
   AOI22_X1 U3388 (.A1(REGISTERS[223]),
	.A2(n2764),
	.B1(REGISTERS[159]),
	.B2(n2763),
	.ZN(n2755));
   AOI22_X1 U3389 (.A1(REGISTERS[127]),
	.A2(FE_OFN8_n2766),
	.B1(REGISTERS[63]),
	.B2(FE_OFN51_n2765),
	.ZN(n2754));
   AOI22_X1 U3390 (.A1(REGISTERS[255]),
	.A2(FE_OFN113_n2768),
	.B1(REGISTERS[191]),
	.B2(FE_OFN11_n2767),
	.ZN(n2753));
   AND4_X1 U3391 (.A1(n2756),
	.A2(n2755),
	.A3(n2754),
	.A4(n2753),
	.ZN(n2779));
   AOI22_X1 U3392 (.A1(REGISTERS[863]),
	.A2(FE_OFN13_n2762),
	.B1(REGISTERS[799]),
	.B2(FE_OFN135_n2761),
	.ZN(n2760));
   AOI22_X1 U3393 (.A1(REGISTERS[991]),
	.A2(FE_OFN54_n2764),
	.B1(REGISTERS[927]),
	.B2(FE_OFN110_n2763),
	.ZN(n2759));
   AOI22_X1 U3394 (.A1(REGISTERS[895]),
	.A2(FE_OFN8_n2766),
	.B1(REGISTERS[831]),
	.B2(FE_OFN51_n2765),
	.ZN(n2758));
   AOI22_X1 U3395 (.A1(REGISTERS[1023]),
	.A2(FE_OFN113_n2768),
	.B1(REGISTERS[959]),
	.B2(FE_OFN11_n2767),
	.ZN(n2757));
   NAND4_X1 U3396 (.A1(n2760),
	.A2(n2759),
	.A3(n2758),
	.A4(n2757),
	.ZN(n2775));
   AOI22_X1 U3397 (.A1(REGISTERS[607]),
	.A2(FE_OFN13_n2762),
	.B1(REGISTERS[543]),
	.B2(FE_OFN135_n2761),
	.ZN(n2772));
   AOI22_X1 U3398 (.A1(REGISTERS[735]),
	.A2(FE_OFN54_n2764),
	.B1(REGISTERS[671]),
	.B2(FE_OFN110_n2763),
	.ZN(n2771));
   AOI22_X1 U3399 (.A1(REGISTERS[639]),
	.A2(FE_OFN8_n2766),
	.B1(REGISTERS[575]),
	.B2(FE_OFN51_n2765),
	.ZN(n2770));
   AOI22_X1 U3400 (.A1(REGISTERS[767]),
	.A2(FE_OFN113_n2768),
	.B1(REGISTERS[703]),
	.B2(FE_OFN11_n2767),
	.ZN(n2769));
   NAND4_X1 U3401 (.A1(n2772),
	.A2(n2771),
	.A3(n2770),
	.A4(n2769),
	.ZN(n2773));
   AOI22_X1 U3402 (.A1(FE_OFN32_n2776),
	.A2(n2775),
	.B1(FE_OFN30_n2774),
	.B2(n2773),
	.ZN(n2777));
   OAI221_X1 U3403 (.A(n2777),
	.B1(n2781),
	.B2(n2780),
	.C1(n2779),
	.C2(n2778),
	.ZN(N31));
   NAND2_X1 U3412 (.A1(ADD_RD2[4]),
	.A2(n3593),
	.ZN(n3588));
   NOR2_X1 U3413 (.A1(n3592),
	.A2(ADD_RD2[1]),
	.ZN(n2902));
   AND2_X2 U3414 (.A1(n2902),
	.A2(ADD_RD2[0]),
	.ZN(n3570));
   NOR2_X1 U3415 (.A1(n3592),
	.A2(n3591),
	.ZN(n2903));
   AND2_X2 U3416 (.A1(ADD_RD2[0]),
	.A2(n2903),
	.ZN(n3569));
   AOI22_X1 U3417 (.A1(REGISTERS[320]),
	.A2(FE_OFN131_n3570),
	.B1(REGISTERS[256]),
	.B2(n3569),
	.ZN(n2909));
   NOR2_X1 U3418 (.A1(ADD_RD2[1]),
	.A2(ADD_RD2[2]),
	.ZN(n2904));
   AND2_X2 U3419 (.A1(n2904),
	.A2(ADD_RD2[0]),
	.ZN(n3572));
   NOR2_X1 U3420 (.A1(n3591),
	.A2(ADD_RD2[2]),
	.ZN(n2905));
   AND2_X2 U3421 (.A1(n2905),
	.A2(ADD_RD2[0]),
	.ZN(n3571));
   AOI22_X1 U3422 (.A1(REGISTERS[448]),
	.A2(FE_OFN46_n3572),
	.B1(REGISTERS[384]),
	.B2(FE_OFN6_n3571),
	.ZN(n2908));
   AND2_X2 U3423 (.A1(n2902),
	.A2(n3590),
	.ZN(n3574));
   AND2_X2 U3424 (.A1(n2903),
	.A2(n3590),
	.ZN(n3573));
   AOI22_X1 U3425 (.A1(REGISTERS[352]),
	.A2(FE_OFN4_n3574),
	.B1(REGISTERS[288]),
	.B2(FE_OFN133_n3573),
	.ZN(n2907));
   AND2_X2 U3426 (.A1(n2904),
	.A2(n3590),
	.ZN(n3576));
   AND2_X2 U3427 (.A1(n2905),
	.A2(n3590),
	.ZN(n3575));
   AOI22_X1 U3428 (.A1(REGISTERS[480]),
	.A2(n3576),
	.B1(REGISTERS[416]),
	.B2(n3575),
	.ZN(n2906));
   AND4_X1 U3429 (.A1(n2909),
	.A2(n2908),
	.A3(n2907),
	.A4(n2906),
	.ZN(n2926));
   NAND2_X2 U3430 (.A1(ADD_RD2[4]),
	.A2(ADD_RD2[3]),
	.ZN(n3586));
   AOI22_X1 U3431 (.A1(REGISTERS[64]),
	.A2(FE_OFN131_n3570),
	.B1(REGISTERS[0]),
	.B2(n3569),
	.ZN(n2913));
   AOI22_X1 U3432 (.A1(REGISTERS[192]),
	.A2(FE_OFN46_n3572),
	.B1(REGISTERS[128]),
	.B2(FE_OFN6_n3571),
	.ZN(n2912));
   AOI22_X1 U3433 (.A1(REGISTERS[96]),
	.A2(FE_OFN4_n3574),
	.B1(REGISTERS[32]),
	.B2(FE_OFN133_n3573),
	.ZN(n2911));
   AOI22_X1 U3434 (.A1(REGISTERS[224]),
	.A2(n3576),
	.B1(REGISTERS[160]),
	.B2(n3575),
	.ZN(n2910));
   AND4_X1 U3435 (.A1(n2913),
	.A2(n2912),
	.A3(n2911),
	.A4(n2910),
	.ZN(n2925));
   AOI22_X1 U3436 (.A1(REGISTERS[832]),
	.A2(n3570),
	.B1(REGISTERS[768]),
	.B2(n3569),
	.ZN(n2917));
   AOI22_X1 U3437 (.A1(REGISTERS[960]),
	.A2(FE_OFN46_n3572),
	.B1(REGISTERS[896]),
	.B2(FE_OFN6_n3571),
	.ZN(n2916));
   AOI22_X1 U3438 (.A1(REGISTERS[864]),
	.A2(FE_OFN4_n3574),
	.B1(REGISTERS[800]),
	.B2(FE_OFN133_n3573),
	.ZN(n2915));
   AOI22_X1 U3439 (.A1(REGISTERS[992]),
	.A2(n3576),
	.B1(REGISTERS[928]),
	.B2(n3575),
	.ZN(n2914));
   NAND4_X1 U3440 (.A1(n2917),
	.A2(n2916),
	.A3(n2915),
	.A4(n2914),
	.ZN(n2923));
   NOR2_X1 U3441 (.A1(ADD_RD2[3]),
	.A2(ADD_RD2[4]),
	.ZN(n3584));
   AOI22_X1 U3442 (.A1(REGISTERS[576]),
	.A2(n3570),
	.B1(REGISTERS[512]),
	.B2(n3569),
	.ZN(n2921));
   AOI22_X1 U3443 (.A1(REGISTERS[704]),
	.A2(FE_OFN46_n3572),
	.B1(REGISTERS[640]),
	.B2(FE_OFN6_n3571),
	.ZN(n2920));
   AOI22_X1 U3444 (.A1(REGISTERS[608]),
	.A2(FE_OFN4_n3574),
	.B1(REGISTERS[544]),
	.B2(FE_OFN133_n3573),
	.ZN(n2919));
   AOI22_X1 U3445 (.A1(REGISTERS[736]),
	.A2(n3576),
	.B1(REGISTERS[672]),
	.B2(n3575),
	.ZN(n2918));
   NAND4_X1 U3446 (.A1(n2921),
	.A2(n2920),
	.A3(n2919),
	.A4(n2918),
	.ZN(n2922));
   NOR2_X1 U3447 (.A1(n3593),
	.A2(ADD_RD2[4]),
	.ZN(n3582));
   AOI22_X1 U3448 (.A1(n2923),
	.A2(FE_OFN33_n3584),
	.B1(n2922),
	.B2(FE_OFN31_n3582),
	.ZN(n2924));
   OAI221_X1 U3449 (.A(n2924),
	.B1(FE_OFN38_n3588),
	.B2(n2926),
	.C1(n3586),
	.C2(n2925),
	.ZN(N127));
   AOI22_X1 U3450 (.A1(REGISTERS[321]),
	.A2(FE_OFN131_n3570),
	.B1(REGISTERS[257]),
	.B2(FE_OFN108_n3569),
	.ZN(n2930));
   AOI22_X1 U3451 (.A1(REGISTERS[449]),
	.A2(n3572),
	.B1(REGISTERS[385]),
	.B2(n3571),
	.ZN(n2929));
   AOI22_X1 U3452 (.A1(REGISTERS[353]),
	.A2(n3574),
	.B1(REGISTERS[289]),
	.B2(n3573),
	.ZN(n2928));
   AOI22_X1 U3453 (.A1(REGISTERS[481]),
	.A2(FE_OFN105_n3576),
	.B1(REGISTERS[417]),
	.B2(FE_OFN48_n3575),
	.ZN(n2927));
   AND4_X1 U3454 (.A1(n2930),
	.A2(n2929),
	.A3(n2928),
	.A4(n2927),
	.ZN(n2947));
   AOI22_X1 U3455 (.A1(REGISTERS[65]),
	.A2(FE_OFN131_n3570),
	.B1(REGISTERS[1]),
	.B2(FE_OFN108_n3569),
	.ZN(n2934));
   AOI22_X1 U3456 (.A1(REGISTERS[193]),
	.A2(n3572),
	.B1(REGISTERS[129]),
	.B2(n3571),
	.ZN(n2933));
   AOI22_X1 U3457 (.A1(REGISTERS[97]),
	.A2(n3574),
	.B1(REGISTERS[33]),
	.B2(n3573),
	.ZN(n2932));
   AOI22_X1 U3458 (.A1(REGISTERS[225]),
	.A2(FE_OFN105_n3576),
	.B1(REGISTERS[161]),
	.B2(FE_OFN48_n3575),
	.ZN(n2931));
   AND4_X1 U3459 (.A1(n2934),
	.A2(n2933),
	.A3(n2932),
	.A4(n2931),
	.ZN(n2946));
   AOI22_X1 U3460 (.A1(REGISTERS[833]),
	.A2(FE_OFN131_n3570),
	.B1(REGISTERS[769]),
	.B2(FE_OFN108_n3569),
	.ZN(n2938));
   AOI22_X1 U3461 (.A1(REGISTERS[961]),
	.A2(FE_OFN46_n3572),
	.B1(REGISTERS[897]),
	.B2(FE_OFN6_n3571),
	.ZN(n2937));
   AOI22_X1 U3462 (.A1(REGISTERS[865]),
	.A2(FE_OFN3_n3574),
	.B1(REGISTERS[801]),
	.B2(FE_OFN133_n3573),
	.ZN(n2936));
   AOI22_X1 U3463 (.A1(REGISTERS[993]),
	.A2(FE_OFN105_n3576),
	.B1(REGISTERS[929]),
	.B2(FE_OFN48_n3575),
	.ZN(n2935));
   NAND4_X1 U3464 (.A1(n2938),
	.A2(n2937),
	.A3(n2936),
	.A4(n2935),
	.ZN(n2944));
   AOI22_X1 U3465 (.A1(REGISTERS[577]),
	.A2(FE_OFN131_n3570),
	.B1(REGISTERS[513]),
	.B2(FE_OFN108_n3569),
	.ZN(n2942));
   AOI22_X1 U3466 (.A1(REGISTERS[705]),
	.A2(FE_OFN46_n3572),
	.B1(REGISTERS[641]),
	.B2(FE_OFN6_n3571),
	.ZN(n2941));
   AOI22_X1 U3467 (.A1(REGISTERS[609]),
	.A2(FE_OFN3_n3574),
	.B1(REGISTERS[545]),
	.B2(FE_OFN133_n3573),
	.ZN(n2940));
   AOI22_X1 U3468 (.A1(REGISTERS[737]),
	.A2(FE_OFN105_n3576),
	.B1(REGISTERS[673]),
	.B2(FE_OFN48_n3575),
	.ZN(n2939));
   NAND4_X1 U3469 (.A1(n2942),
	.A2(n2941),
	.A3(n2940),
	.A4(n2939),
	.ZN(n2943));
   AOI22_X1 U3470 (.A1(n2944),
	.A2(FE_OFN33_n3584),
	.B1(n2943),
	.B2(FE_OFN31_n3582),
	.ZN(n2945));
   OAI221_X1 U3471 (.A(n2945),
	.B1(FE_OFN38_n3588),
	.B2(n2947),
	.C1(n3586),
	.C2(n2946),
	.ZN(N126));
   AOI22_X1 U3472 (.A1(REGISTERS[322]),
	.A2(FE_OFN131_n3570),
	.B1(REGISTERS[258]),
	.B2(n3569),
	.ZN(n2951));
   AOI22_X1 U3473 (.A1(REGISTERS[450]),
	.A2(FE_OFN46_n3572),
	.B1(REGISTERS[386]),
	.B2(FE_OFN6_n3571),
	.ZN(n2950));
   AOI22_X1 U3474 (.A1(REGISTERS[354]),
	.A2(FE_OFN4_n3574),
	.B1(REGISTERS[290]),
	.B2(FE_OFN134_n3573),
	.ZN(n2949));
   AOI22_X1 U3475 (.A1(REGISTERS[482]),
	.A2(FE_OFN105_n3576),
	.B1(REGISTERS[418]),
	.B2(FE_OFN48_n3575),
	.ZN(n2948));
   AND4_X1 U3476 (.A1(n2951),
	.A2(n2950),
	.A3(n2949),
	.A4(n2948),
	.ZN(n2968));
   AOI22_X1 U3477 (.A1(REGISTERS[66]),
	.A2(FE_OFN131_n3570),
	.B1(REGISTERS[2]),
	.B2(n3569),
	.ZN(n2955));
   AOI22_X1 U3478 (.A1(REGISTERS[194]),
	.A2(FE_OFN46_n3572),
	.B1(REGISTERS[130]),
	.B2(FE_OFN6_n3571),
	.ZN(n2954));
   AOI22_X1 U3479 (.A1(REGISTERS[98]),
	.A2(FE_OFN4_n3574),
	.B1(REGISTERS[34]),
	.B2(FE_OFN134_n3573),
	.ZN(n2953));
   AOI22_X1 U3480 (.A1(REGISTERS[226]),
	.A2(FE_OFN105_n3576),
	.B1(REGISTERS[162]),
	.B2(FE_OFN48_n3575),
	.ZN(n2952));
   AND4_X1 U3481 (.A1(n2955),
	.A2(n2954),
	.A3(n2953),
	.A4(n2952),
	.ZN(n2967));
   AOI22_X1 U3482 (.A1(REGISTERS[834]),
	.A2(FE_OFN132_n3570),
	.B1(REGISTERS[770]),
	.B2(FE_OFN109_n3569),
	.ZN(n2959));
   AOI22_X1 U3483 (.A1(REGISTERS[962]),
	.A2(FE_OFN47_n3572),
	.B1(REGISTERS[898]),
	.B2(FE_OFN7_n3571),
	.ZN(n2958));
   AOI22_X1 U3484 (.A1(REGISTERS[866]),
	.A2(FE_OFN5_n3574),
	.B1(REGISTERS[802]),
	.B2(FE_OFN134_n3573),
	.ZN(n2957));
   AOI22_X1 U3485 (.A1(REGISTERS[994]),
	.A2(FE_OFN107_n3576),
	.B1(REGISTERS[930]),
	.B2(FE_OFN49_n3575),
	.ZN(n2956));
   NAND4_X1 U3486 (.A1(n2959),
	.A2(n2958),
	.A3(n2957),
	.A4(n2956),
	.ZN(n2965));
   AOI22_X1 U3487 (.A1(REGISTERS[578]),
	.A2(FE_OFN132_n3570),
	.B1(REGISTERS[514]),
	.B2(FE_OFN109_n3569),
	.ZN(n2963));
   AOI22_X1 U3488 (.A1(REGISTERS[706]),
	.A2(FE_OFN47_n3572),
	.B1(REGISTERS[642]),
	.B2(FE_OFN7_n3571),
	.ZN(n2962));
   AOI22_X1 U3489 (.A1(REGISTERS[610]),
	.A2(FE_OFN5_n3574),
	.B1(REGISTERS[546]),
	.B2(FE_OFN134_n3573),
	.ZN(n2961));
   AOI22_X1 U3490 (.A1(REGISTERS[738]),
	.A2(FE_OFN107_n3576),
	.B1(REGISTERS[674]),
	.B2(FE_OFN49_n3575),
	.ZN(n2960));
   NAND4_X1 U3491 (.A1(n2963),
	.A2(n2962),
	.A3(n2961),
	.A4(n2960),
	.ZN(n2964));
   AOI22_X1 U3492 (.A1(n2965),
	.A2(FE_OFN33_n3584),
	.B1(n2964),
	.B2(FE_OFN31_n3582),
	.ZN(n2966));
   OAI221_X1 U3493 (.A(n2966),
	.B1(FE_OFN38_n3588),
	.B2(n2968),
	.C1(n3586),
	.C2(n2967),
	.ZN(N125));
   AOI22_X1 U3494 (.A1(REGISTERS[323]),
	.A2(FE_OFN132_n3570),
	.B1(REGISTERS[259]),
	.B2(FE_OFN109_n3569),
	.ZN(n2972));
   AOI22_X1 U3495 (.A1(REGISTERS[451]),
	.A2(FE_OFN47_n3572),
	.B1(REGISTERS[387]),
	.B2(FE_OFN6_n3571),
	.ZN(n2971));
   AOI22_X1 U3496 (.A1(REGISTERS[355]),
	.A2(FE_OFN4_n3574),
	.B1(REGISTERS[291]),
	.B2(FE_OFN133_n3573),
	.ZN(n2970));
   AOI22_X1 U3497 (.A1(REGISTERS[483]),
	.A2(FE_OFN107_n3576),
	.B1(REGISTERS[419]),
	.B2(FE_OFN50_n3575),
	.ZN(n2969));
   AND4_X1 U3498 (.A1(n2972),
	.A2(n2971),
	.A3(n2970),
	.A4(n2969),
	.ZN(n2989));
   AOI22_X1 U3499 (.A1(REGISTERS[67]),
	.A2(FE_OFN132_n3570),
	.B1(REGISTERS[3]),
	.B2(FE_OFN109_n3569),
	.ZN(n2976));
   AOI22_X1 U3500 (.A1(REGISTERS[195]),
	.A2(FE_OFN47_n3572),
	.B1(REGISTERS[131]),
	.B2(FE_OFN6_n3571),
	.ZN(n2975));
   AOI22_X1 U3501 (.A1(REGISTERS[99]),
	.A2(FE_OFN4_n3574),
	.B1(REGISTERS[35]),
	.B2(FE_OFN134_n3573),
	.ZN(n2974));
   AOI22_X1 U3502 (.A1(REGISTERS[227]),
	.A2(FE_OFN107_n3576),
	.B1(REGISTERS[163]),
	.B2(FE_OFN50_n3575),
	.ZN(n2973));
   AND4_X1 U3503 (.A1(n2976),
	.A2(n2975),
	.A3(n2974),
	.A4(n2973),
	.ZN(n2988));
   AOI22_X1 U3504 (.A1(REGISTERS[835]),
	.A2(FE_OFN132_n3570),
	.B1(REGISTERS[771]),
	.B2(FE_OFN109_n3569),
	.ZN(n2980));
   AOI22_X1 U3505 (.A1(REGISTERS[963]),
	.A2(FE_OFN47_n3572),
	.B1(REGISTERS[899]),
	.B2(FE_OFN7_n3571),
	.ZN(n2979));
   AOI22_X1 U3506 (.A1(REGISTERS[867]),
	.A2(FE_OFN5_n3574),
	.B1(REGISTERS[803]),
	.B2(FE_OFN134_n3573),
	.ZN(n2978));
   AOI22_X1 U3507 (.A1(REGISTERS[995]),
	.A2(FE_OFN107_n3576),
	.B1(REGISTERS[931]),
	.B2(FE_OFN49_n3575),
	.ZN(n2977));
   NAND4_X1 U3508 (.A1(n2980),
	.A2(n2979),
	.A3(n2978),
	.A4(n2977),
	.ZN(n2986));
   AOI22_X1 U3509 (.A1(REGISTERS[579]),
	.A2(FE_OFN132_n3570),
	.B1(REGISTERS[515]),
	.B2(FE_OFN109_n3569),
	.ZN(n2984));
   AOI22_X1 U3510 (.A1(REGISTERS[707]),
	.A2(FE_OFN47_n3572),
	.B1(REGISTERS[643]),
	.B2(FE_OFN7_n3571),
	.ZN(n2983));
   AOI22_X1 U3511 (.A1(REGISTERS[611]),
	.A2(FE_OFN5_n3574),
	.B1(REGISTERS[547]),
	.B2(FE_OFN134_n3573),
	.ZN(n2982));
   AOI22_X1 U3512 (.A1(REGISTERS[739]),
	.A2(FE_OFN107_n3576),
	.B1(REGISTERS[675]),
	.B2(FE_OFN49_n3575),
	.ZN(n2981));
   NAND4_X1 U3513 (.A1(n2984),
	.A2(n2983),
	.A3(n2982),
	.A4(n2981),
	.ZN(n2985));
   AOI22_X1 U3514 (.A1(n2986),
	.A2(FE_OFN33_n3584),
	.B1(n2985),
	.B2(FE_OFN31_n3582),
	.ZN(n2987));
   OAI221_X1 U3515 (.A(n2987),
	.B1(FE_OFN38_n3588),
	.B2(n2989),
	.C1(n3586),
	.C2(n2988),
	.ZN(N124));
   AOI22_X1 U3516 (.A1(REGISTERS[324]),
	.A2(n3570),
	.B1(REGISTERS[260]),
	.B2(n3569),
	.ZN(n2993));
   AOI22_X1 U3517 (.A1(REGISTERS[452]),
	.A2(n3572),
	.B1(REGISTERS[388]),
	.B2(n3571),
	.ZN(n2992));
   AOI22_X1 U3518 (.A1(REGISTERS[356]),
	.A2(n3574),
	.B1(REGISTERS[292]),
	.B2(n3573),
	.ZN(n2991));
   AOI22_X1 U3519 (.A1(REGISTERS[484]),
	.A2(n3576),
	.B1(REGISTERS[420]),
	.B2(n3575),
	.ZN(n2990));
   AND4_X1 U3520 (.A1(n2993),
	.A2(n2992),
	.A3(n2991),
	.A4(n2990),
	.ZN(n3010));
   AOI22_X1 U3521 (.A1(REGISTERS[68]),
	.A2(n3570),
	.B1(REGISTERS[4]),
	.B2(FE_OFN108_n3569),
	.ZN(n2997));
   AOI22_X1 U3522 (.A1(REGISTERS[196]),
	.A2(n3572),
	.B1(REGISTERS[132]),
	.B2(n3571),
	.ZN(n2996));
   AOI22_X1 U3523 (.A1(REGISTERS[100]),
	.A2(n3574),
	.B1(REGISTERS[36]),
	.B2(n3573),
	.ZN(n2995));
   AOI22_X1 U3524 (.A1(REGISTERS[228]),
	.A2(n3576),
	.B1(REGISTERS[164]),
	.B2(n3575),
	.ZN(n2994));
   AND4_X1 U3525 (.A1(n2997),
	.A2(n2996),
	.A3(n2995),
	.A4(n2994),
	.ZN(n3009));
   AOI22_X1 U3526 (.A1(REGISTERS[836]),
	.A2(n3570),
	.B1(REGISTERS[772]),
	.B2(n3569),
	.ZN(n3001));
   AOI22_X1 U3527 (.A1(REGISTERS[964]),
	.A2(FE_OFN46_n3572),
	.B1(REGISTERS[900]),
	.B2(FE_OFN6_n3571),
	.ZN(n3000));
   AOI22_X1 U3528 (.A1(REGISTERS[868]),
	.A2(FE_OFN4_n3574),
	.B1(REGISTERS[804]),
	.B2(n3573),
	.ZN(n2999));
   AOI22_X1 U3529 (.A1(REGISTERS[996]),
	.A2(n3576),
	.B1(REGISTERS[932]),
	.B2(n3575),
	.ZN(n2998));
   NAND4_X1 U3530 (.A1(n3001),
	.A2(n3000),
	.A3(n2999),
	.A4(n2998),
	.ZN(n3007));
   AOI22_X1 U3531 (.A1(REGISTERS[580]),
	.A2(n3570),
	.B1(REGISTERS[516]),
	.B2(n3569),
	.ZN(n3005));
   AOI22_X1 U3532 (.A1(REGISTERS[708]),
	.A2(FE_OFN46_n3572),
	.B1(REGISTERS[644]),
	.B2(FE_OFN6_n3571),
	.ZN(n3004));
   AOI22_X1 U3533 (.A1(REGISTERS[612]),
	.A2(FE_OFN4_n3574),
	.B1(REGISTERS[548]),
	.B2(FE_OFN133_n3573),
	.ZN(n3003));
   AOI22_X1 U3534 (.A1(REGISTERS[740]),
	.A2(n3576),
	.B1(REGISTERS[676]),
	.B2(n3575),
	.ZN(n3002));
   NAND4_X1 U3535 (.A1(n3005),
	.A2(n3004),
	.A3(n3003),
	.A4(n3002),
	.ZN(n3006));
   AOI22_X1 U3536 (.A1(n3007),
	.A2(FE_OFN33_n3584),
	.B1(n3006),
	.B2(FE_OFN31_n3582),
	.ZN(n3008));
   OAI221_X1 U3537 (.A(n3008),
	.B1(FE_OFN38_n3588),
	.B2(n3010),
	.C1(n3586),
	.C2(n3009),
	.ZN(N123));
   AOI22_X1 U3538 (.A1(REGISTERS[325]),
	.A2(FE_OFN132_n3570),
	.B1(REGISTERS[261]),
	.B2(FE_OFN109_n3569),
	.ZN(n3014));
   AOI22_X1 U3539 (.A1(REGISTERS[453]),
	.A2(FE_OFN47_n3572),
	.B1(REGISTERS[389]),
	.B2(FE_OFN6_n3571),
	.ZN(n3013));
   AOI22_X1 U3540 (.A1(REGISTERS[357]),
	.A2(FE_OFN4_n3574),
	.B1(REGISTERS[293]),
	.B2(FE_OFN133_n3573),
	.ZN(n3012));
   AOI22_X1 U3541 (.A1(REGISTERS[485]),
	.A2(FE_OFN107_n3576),
	.B1(REGISTERS[421]),
	.B2(FE_OFN50_n3575),
	.ZN(n3011));
   AND4_X1 U3542 (.A1(n3014),
	.A2(n3013),
	.A3(n3012),
	.A4(n3011),
	.ZN(n3031));
   AOI22_X1 U3543 (.A1(REGISTERS[69]),
	.A2(FE_OFN132_n3570),
	.B1(REGISTERS[5]),
	.B2(FE_OFN109_n3569),
	.ZN(n3018));
   AOI22_X1 U3544 (.A1(REGISTERS[197]),
	.A2(FE_OFN47_n3572),
	.B1(REGISTERS[133]),
	.B2(FE_OFN6_n3571),
	.ZN(n3017));
   AOI22_X1 U3545 (.A1(REGISTERS[101]),
	.A2(FE_OFN4_n3574),
	.B1(REGISTERS[37]),
	.B2(FE_OFN133_n3573),
	.ZN(n3016));
   AOI22_X1 U3546 (.A1(REGISTERS[229]),
	.A2(FE_OFN107_n3576),
	.B1(REGISTERS[165]),
	.B2(FE_OFN50_n3575),
	.ZN(n3015));
   AND4_X1 U3547 (.A1(n3018),
	.A2(n3017),
	.A3(n3016),
	.A4(n3015),
	.ZN(n3030));
   AOI22_X1 U3548 (.A1(REGISTERS[837]),
	.A2(n3570),
	.B1(REGISTERS[773]),
	.B2(n3569),
	.ZN(n3022));
   AOI22_X1 U3549 (.A1(REGISTERS[965]),
	.A2(FE_OFN47_n3572),
	.B1(REGISTERS[901]),
	.B2(FE_OFN7_n3571),
	.ZN(n3021));
   AOI22_X1 U3550 (.A1(REGISTERS[869]),
	.A2(FE_OFN5_n3574),
	.B1(REGISTERS[805]),
	.B2(FE_OFN134_n3573),
	.ZN(n3020));
   AOI22_X1 U3551 (.A1(REGISTERS[997]),
	.A2(FE_OFN107_n3576),
	.B1(REGISTERS[933]),
	.B2(FE_OFN50_n3575),
	.ZN(n3019));
   NAND4_X1 U3552 (.A1(n3022),
	.A2(n3021),
	.A3(n3020),
	.A4(n3019),
	.ZN(n3028));
   AOI22_X1 U3553 (.A1(REGISTERS[581]),
	.A2(n3570),
	.B1(REGISTERS[517]),
	.B2(n3569),
	.ZN(n3026));
   AOI22_X1 U3554 (.A1(REGISTERS[709]),
	.A2(FE_OFN47_n3572),
	.B1(REGISTERS[645]),
	.B2(FE_OFN7_n3571),
	.ZN(n3025));
   AOI22_X1 U3555 (.A1(REGISTERS[613]),
	.A2(FE_OFN5_n3574),
	.B1(REGISTERS[549]),
	.B2(FE_OFN134_n3573),
	.ZN(n3024));
   AOI22_X1 U3556 (.A1(REGISTERS[741]),
	.A2(FE_OFN107_n3576),
	.B1(REGISTERS[677]),
	.B2(FE_OFN50_n3575),
	.ZN(n3023));
   NAND4_X1 U3557 (.A1(n3026),
	.A2(n3025),
	.A3(n3024),
	.A4(n3023),
	.ZN(n3027));
   AOI22_X1 U3558 (.A1(n3028),
	.A2(FE_OFN33_n3584),
	.B1(n3027),
	.B2(FE_OFN31_n3582),
	.ZN(n3029));
   OAI221_X1 U3559 (.A(n3029),
	.B1(FE_OFN38_n3588),
	.B2(n3031),
	.C1(n3586),
	.C2(n3030),
	.ZN(N122));
   AOI22_X1 U3560 (.A1(REGISTERS[326]),
	.A2(FE_OFN131_n3570),
	.B1(REGISTERS[262]),
	.B2(FE_OFN108_n3569),
	.ZN(n3035));
   AOI22_X1 U3561 (.A1(REGISTERS[454]),
	.A2(n3572),
	.B1(REGISTERS[390]),
	.B2(n3571),
	.ZN(n3034));
   AOI22_X1 U3562 (.A1(REGISTERS[358]),
	.A2(n3574),
	.B1(REGISTERS[294]),
	.B2(n3573),
	.ZN(n3033));
   AOI22_X1 U3563 (.A1(REGISTERS[486]),
	.A2(n3576),
	.B1(REGISTERS[422]),
	.B2(FE_OFN48_n3575),
	.ZN(n3032));
   AND4_X1 U3564 (.A1(n3035),
	.A2(n3034),
	.A3(n3033),
	.A4(n3032),
	.ZN(n3052));
   AOI22_X1 U3565 (.A1(REGISTERS[70]),
	.A2(FE_OFN131_n3570),
	.B1(REGISTERS[6]),
	.B2(FE_OFN108_n3569),
	.ZN(n3039));
   AOI22_X1 U3566 (.A1(REGISTERS[198]),
	.A2(n3572),
	.B1(REGISTERS[134]),
	.B2(n3571),
	.ZN(n3038));
   AOI22_X1 U3567 (.A1(REGISTERS[102]),
	.A2(n3574),
	.B1(REGISTERS[38]),
	.B2(n3573),
	.ZN(n3037));
   AOI22_X1 U3568 (.A1(REGISTERS[230]),
	.A2(FE_OFN105_n3576),
	.B1(REGISTERS[166]),
	.B2(FE_OFN48_n3575),
	.ZN(n3036));
   AND4_X1 U3569 (.A1(n3039),
	.A2(n3038),
	.A3(n3037),
	.A4(n3036),
	.ZN(n3051));
   AOI22_X1 U3570 (.A1(REGISTERS[838]),
	.A2(FE_OFN131_n3570),
	.B1(REGISTERS[774]),
	.B2(FE_OFN108_n3569),
	.ZN(n3043));
   AOI22_X1 U3571 (.A1(REGISTERS[966]),
	.A2(FE_OFN46_n3572),
	.B1(REGISTERS[902]),
	.B2(FE_OFN6_n3571),
	.ZN(n3042));
   AOI22_X1 U3572 (.A1(REGISTERS[870]),
	.A2(FE_OFN3_n3574),
	.B1(REGISTERS[806]),
	.B2(FE_OFN133_n3573),
	.ZN(n3041));
   AOI22_X1 U3573 (.A1(REGISTERS[998]),
	.A2(FE_OFN105_n3576),
	.B1(REGISTERS[934]),
	.B2(FE_OFN48_n3575),
	.ZN(n3040));
   NAND4_X1 U3574 (.A1(n3043),
	.A2(n3042),
	.A3(n3041),
	.A4(n3040),
	.ZN(n3049));
   AOI22_X1 U3575 (.A1(REGISTERS[582]),
	.A2(FE_OFN131_n3570),
	.B1(REGISTERS[518]),
	.B2(n3569),
	.ZN(n3047));
   AOI22_X1 U3576 (.A1(REGISTERS[710]),
	.A2(FE_OFN46_n3572),
	.B1(REGISTERS[646]),
	.B2(FE_OFN6_n3571),
	.ZN(n3046));
   AOI22_X1 U3577 (.A1(REGISTERS[614]),
	.A2(FE_OFN4_n3574),
	.B1(REGISTERS[550]),
	.B2(FE_OFN134_n3573),
	.ZN(n3045));
   AOI22_X1 U3578 (.A1(REGISTERS[742]),
	.A2(FE_OFN105_n3576),
	.B1(REGISTERS[678]),
	.B2(FE_OFN48_n3575),
	.ZN(n3044));
   NAND4_X1 U3579 (.A1(n3047),
	.A2(n3046),
	.A3(n3045),
	.A4(n3044),
	.ZN(n3048));
   AOI22_X1 U3580 (.A1(n3049),
	.A2(FE_OFN33_n3584),
	.B1(n3048),
	.B2(FE_OFN31_n3582),
	.ZN(n3050));
   OAI221_X1 U3581 (.A(n3050),
	.B1(FE_OFN38_n3588),
	.B2(n3052),
	.C1(n3586),
	.C2(n3051),
	.ZN(N121));
   AOI22_X1 U3582 (.A1(REGISTERS[327]),
	.A2(FE_OFN132_n3570),
	.B1(REGISTERS[263]),
	.B2(FE_OFN109_n3569),
	.ZN(n3056));
   AOI22_X1 U3583 (.A1(REGISTERS[455]),
	.A2(FE_OFN47_n3572),
	.B1(REGISTERS[391]),
	.B2(FE_OFN6_n3571),
	.ZN(n3055));
   AOI22_X1 U3584 (.A1(REGISTERS[359]),
	.A2(FE_OFN4_n3574),
	.B1(REGISTERS[295]),
	.B2(FE_OFN133_n3573),
	.ZN(n3054));
   AOI22_X1 U3585 (.A1(REGISTERS[487]),
	.A2(FE_OFN107_n3576),
	.B1(REGISTERS[423]),
	.B2(FE_OFN50_n3575),
	.ZN(n3053));
   AND4_X1 U3586 (.A1(n3056),
	.A2(n3055),
	.A3(n3054),
	.A4(n3053),
	.ZN(n3073));
   AOI22_X1 U3587 (.A1(REGISTERS[71]),
	.A2(FE_OFN132_n3570),
	.B1(REGISTERS[7]),
	.B2(FE_OFN109_n3569),
	.ZN(n3060));
   AOI22_X1 U3588 (.A1(REGISTERS[199]),
	.A2(FE_OFN47_n3572),
	.B1(REGISTERS[135]),
	.B2(FE_OFN6_n3571),
	.ZN(n3059));
   AOI22_X1 U3589 (.A1(REGISTERS[103]),
	.A2(FE_OFN4_n3574),
	.B1(REGISTERS[39]),
	.B2(FE_OFN133_n3573),
	.ZN(n3058));
   AOI22_X1 U3590 (.A1(REGISTERS[231]),
	.A2(FE_OFN107_n3576),
	.B1(REGISTERS[167]),
	.B2(FE_OFN50_n3575),
	.ZN(n3057));
   AND4_X1 U3591 (.A1(n3060),
	.A2(n3059),
	.A3(n3058),
	.A4(n3057),
	.ZN(n3072));
   AOI22_X1 U3592 (.A1(REGISTERS[839]),
	.A2(FE_OFN132_n3570),
	.B1(REGISTERS[775]),
	.B2(FE_OFN109_n3569),
	.ZN(n3064));
   AOI22_X1 U3593 (.A1(REGISTERS[967]),
	.A2(FE_OFN47_n3572),
	.B1(REGISTERS[903]),
	.B2(FE_OFN7_n3571),
	.ZN(n3063));
   AOI22_X1 U3594 (.A1(REGISTERS[871]),
	.A2(FE_OFN5_n3574),
	.B1(REGISTERS[807]),
	.B2(FE_OFN134_n3573),
	.ZN(n3062));
   AOI22_X1 U3595 (.A1(REGISTERS[999]),
	.A2(FE_OFN107_n3576),
	.B1(REGISTERS[935]),
	.B2(FE_OFN49_n3575),
	.ZN(n3061));
   NAND4_X1 U3596 (.A1(n3064),
	.A2(n3063),
	.A3(n3062),
	.A4(n3061),
	.ZN(n3070));
   AOI22_X1 U3597 (.A1(REGISTERS[583]),
	.A2(FE_OFN132_n3570),
	.B1(REGISTERS[519]),
	.B2(FE_OFN109_n3569),
	.ZN(n3068));
   AOI22_X1 U3598 (.A1(REGISTERS[711]),
	.A2(FE_OFN47_n3572),
	.B1(REGISTERS[647]),
	.B2(FE_OFN7_n3571),
	.ZN(n3067));
   AOI22_X1 U3599 (.A1(REGISTERS[615]),
	.A2(FE_OFN5_n3574),
	.B1(REGISTERS[551]),
	.B2(FE_OFN134_n3573),
	.ZN(n3066));
   AOI22_X1 U3600 (.A1(REGISTERS[743]),
	.A2(FE_OFN107_n3576),
	.B1(REGISTERS[679]),
	.B2(FE_OFN49_n3575),
	.ZN(n3065));
   NAND4_X1 U3601 (.A1(n3068),
	.A2(n3067),
	.A3(n3066),
	.A4(n3065),
	.ZN(n3069));
   AOI22_X1 U3602 (.A1(n3070),
	.A2(FE_OFN33_n3584),
	.B1(n3069),
	.B2(FE_OFN31_n3582),
	.ZN(n3071));
   OAI221_X1 U3603 (.A(n3071),
	.B1(FE_OFN38_n3588),
	.B2(n3073),
	.C1(n3586),
	.C2(n3072),
	.ZN(N120));
   AOI22_X1 U3604 (.A1(REGISTERS[328]),
	.A2(FE_OFN131_n3570),
	.B1(REGISTERS[264]),
	.B2(FE_OFN108_n3569),
	.ZN(n3077));
   AOI22_X1 U3605 (.A1(REGISTERS[456]),
	.A2(n3572),
	.B1(REGISTERS[392]),
	.B2(n3571),
	.ZN(n3076));
   AOI22_X1 U3606 (.A1(REGISTERS[360]),
	.A2(n3574),
	.B1(REGISTERS[296]),
	.B2(n3573),
	.ZN(n3075));
   AOI22_X1 U3607 (.A1(REGISTERS[488]),
	.A2(n3576),
	.B1(REGISTERS[424]),
	.B2(FE_OFN48_n3575),
	.ZN(n3074));
   AND4_X1 U3608 (.A1(n3077),
	.A2(n3076),
	.A3(n3075),
	.A4(n3074),
	.ZN(n3094));
   AOI22_X1 U3609 (.A1(REGISTERS[72]),
	.A2(FE_OFN131_n3570),
	.B1(REGISTERS[8]),
	.B2(FE_OFN108_n3569),
	.ZN(n3081));
   AOI22_X1 U3610 (.A1(REGISTERS[200]),
	.A2(n3572),
	.B1(REGISTERS[136]),
	.B2(n3571),
	.ZN(n3080));
   AOI22_X1 U3611 (.A1(REGISTERS[104]),
	.A2(n3574),
	.B1(REGISTERS[40]),
	.B2(n3573),
	.ZN(n3079));
   AOI22_X1 U3612 (.A1(REGISTERS[232]),
	.A2(n3576),
	.B1(REGISTERS[168]),
	.B2(FE_OFN48_n3575),
	.ZN(n3078));
   AND4_X1 U3613 (.A1(n3081),
	.A2(n3080),
	.A3(n3079),
	.A4(n3078),
	.ZN(n3093));
   AOI22_X1 U3614 (.A1(REGISTERS[840]),
	.A2(FE_OFN131_n3570),
	.B1(REGISTERS[776]),
	.B2(FE_OFN108_n3569),
	.ZN(n3085));
   AOI22_X1 U3615 (.A1(REGISTERS[968]),
	.A2(FE_OFN46_n3572),
	.B1(REGISTERS[904]),
	.B2(FE_OFN6_n3571),
	.ZN(n3084));
   AOI22_X1 U3616 (.A1(REGISTERS[872]),
	.A2(FE_OFN3_n3574),
	.B1(REGISTERS[808]),
	.B2(FE_OFN133_n3573),
	.ZN(n3083));
   AOI22_X1 U3617 (.A1(REGISTERS[1000]),
	.A2(n3576),
	.B1(REGISTERS[936]),
	.B2(n3575),
	.ZN(n3082));
   NAND4_X1 U3618 (.A1(n3085),
	.A2(n3084),
	.A3(n3083),
	.A4(n3082),
	.ZN(n3091));
   AOI22_X1 U3619 (.A1(REGISTERS[584]),
	.A2(FE_OFN131_n3570),
	.B1(REGISTERS[520]),
	.B2(FE_OFN108_n3569),
	.ZN(n3089));
   AOI22_X1 U3620 (.A1(REGISTERS[712]),
	.A2(FE_OFN46_n3572),
	.B1(REGISTERS[648]),
	.B2(FE_OFN6_n3571),
	.ZN(n3088));
   AOI22_X1 U3621 (.A1(REGISTERS[616]),
	.A2(FE_OFN3_n3574),
	.B1(REGISTERS[552]),
	.B2(FE_OFN133_n3573),
	.ZN(n3087));
   AOI22_X1 U3622 (.A1(REGISTERS[744]),
	.A2(n3576),
	.B1(REGISTERS[680]),
	.B2(n3575),
	.ZN(n3086));
   NAND4_X1 U3623 (.A1(n3089),
	.A2(n3088),
	.A3(n3087),
	.A4(n3086),
	.ZN(n3090));
   AOI22_X1 U3624 (.A1(n3091),
	.A2(FE_OFN33_n3584),
	.B1(n3090),
	.B2(FE_OFN31_n3582),
	.ZN(n3092));
   OAI221_X1 U3625 (.A(n3092),
	.B1(FE_OFN38_n3588),
	.B2(n3094),
	.C1(n3586),
	.C2(n3093),
	.ZN(N119));
   AOI22_X1 U3626 (.A1(REGISTERS[329]),
	.A2(n3570),
	.B1(REGISTERS[265]),
	.B2(n3569),
	.ZN(n3098));
   AOI22_X1 U3627 (.A1(REGISTERS[457]),
	.A2(FE_OFN46_n3572),
	.B1(REGISTERS[393]),
	.B2(FE_OFN6_n3571),
	.ZN(n3097));
   AOI22_X1 U3628 (.A1(REGISTERS[361]),
	.A2(FE_OFN4_n3574),
	.B1(REGISTERS[297]),
	.B2(FE_OFN133_n3573),
	.ZN(n3096));
   AOI22_X1 U3629 (.A1(REGISTERS[489]),
	.A2(n3576),
	.B1(REGISTERS[425]),
	.B2(n3575),
	.ZN(n3095));
   AND4_X1 U3630 (.A1(n3098),
	.A2(n3097),
	.A3(n3096),
	.A4(n3095),
	.ZN(n3115));
   AOI22_X1 U3631 (.A1(REGISTERS[73]),
	.A2(n3570),
	.B1(REGISTERS[9]),
	.B2(n3569),
	.ZN(n3102));
   AOI22_X1 U3632 (.A1(REGISTERS[201]),
	.A2(FE_OFN46_n3572),
	.B1(REGISTERS[137]),
	.B2(FE_OFN6_n3571),
	.ZN(n3101));
   AOI22_X1 U3633 (.A1(REGISTERS[105]),
	.A2(FE_OFN4_n3574),
	.B1(REGISTERS[41]),
	.B2(FE_OFN133_n3573),
	.ZN(n3100));
   AOI22_X1 U3634 (.A1(REGISTERS[233]),
	.A2(n3576),
	.B1(REGISTERS[169]),
	.B2(n3575),
	.ZN(n3099));
   AND4_X1 U3635 (.A1(n3102),
	.A2(n3101),
	.A3(n3100),
	.A4(n3099),
	.ZN(n3114));
   AOI22_X1 U3636 (.A1(REGISTERS[841]),
	.A2(n3570),
	.B1(REGISTERS[777]),
	.B2(n3569),
	.ZN(n3106));
   AOI22_X1 U3637 (.A1(REGISTERS[969]),
	.A2(FE_OFN47_n3572),
	.B1(REGISTERS[905]),
	.B2(FE_OFN6_n3571),
	.ZN(n3105));
   AOI22_X1 U3638 (.A1(REGISTERS[873]),
	.A2(FE_OFN4_n3574),
	.B1(REGISTERS[809]),
	.B2(FE_OFN133_n3573),
	.ZN(n3104));
   AOI22_X1 U3639 (.A1(REGISTERS[1001]),
	.A2(n3576),
	.B1(REGISTERS[937]),
	.B2(n3575),
	.ZN(n3103));
   NAND4_X1 U3640 (.A1(n3106),
	.A2(n3105),
	.A3(n3104),
	.A4(n3103),
	.ZN(n3112));
   AOI22_X1 U3641 (.A1(REGISTERS[585]),
	.A2(n3570),
	.B1(REGISTERS[521]),
	.B2(n3569),
	.ZN(n3110));
   AOI22_X1 U3642 (.A1(REGISTERS[713]),
	.A2(FE_OFN46_n3572),
	.B1(REGISTERS[649]),
	.B2(FE_OFN6_n3571),
	.ZN(n3109));
   AOI22_X1 U3643 (.A1(REGISTERS[617]),
	.A2(FE_OFN4_n3574),
	.B1(REGISTERS[553]),
	.B2(FE_OFN133_n3573),
	.ZN(n3108));
   AOI22_X1 U3644 (.A1(REGISTERS[745]),
	.A2(n3576),
	.B1(REGISTERS[681]),
	.B2(n3575),
	.ZN(n3107));
   NAND4_X1 U3645 (.A1(n3110),
	.A2(n3109),
	.A3(n3108),
	.A4(n3107),
	.ZN(n3111));
   AOI22_X1 U3646 (.A1(n3112),
	.A2(FE_OFN33_n3584),
	.B1(n3111),
	.B2(FE_OFN31_n3582),
	.ZN(n3113));
   OAI221_X1 U3647 (.A(n3113),
	.B1(FE_OFN38_n3588),
	.B2(n3115),
	.C1(n3586),
	.C2(n3114),
	.ZN(N118));
   AOI22_X1 U3648 (.A1(REGISTERS[330]),
	.A2(n3570),
	.B1(REGISTERS[266]),
	.B2(FE_OFN108_n3569),
	.ZN(n3119));
   AOI22_X1 U3649 (.A1(REGISTERS[458]),
	.A2(n3572),
	.B1(REGISTERS[394]),
	.B2(n3571),
	.ZN(n3118));
   AOI22_X1 U3650 (.A1(REGISTERS[362]),
	.A2(n3574),
	.B1(REGISTERS[298]),
	.B2(n3573),
	.ZN(n3117));
   AOI22_X1 U3651 (.A1(REGISTERS[490]),
	.A2(n3576),
	.B1(REGISTERS[426]),
	.B2(n3575),
	.ZN(n3116));
   AND4_X1 U3652 (.A1(n3119),
	.A2(n3118),
	.A3(n3117),
	.A4(n3116),
	.ZN(n3136));
   AOI22_X1 U3653 (.A1(REGISTERS[74]),
	.A2(n3570),
	.B1(REGISTERS[10]),
	.B2(FE_OFN108_n3569),
	.ZN(n3123));
   AOI22_X1 U3654 (.A1(REGISTERS[202]),
	.A2(n3572),
	.B1(REGISTERS[138]),
	.B2(n3571),
	.ZN(n3122));
   AOI22_X1 U3655 (.A1(REGISTERS[106]),
	.A2(n3574),
	.B1(REGISTERS[42]),
	.B2(n3573),
	.ZN(n3121));
   AOI22_X1 U3656 (.A1(REGISTERS[234]),
	.A2(n3576),
	.B1(REGISTERS[170]),
	.B2(n3575),
	.ZN(n3120));
   AND4_X1 U3657 (.A1(n3123),
	.A2(n3122),
	.A3(n3121),
	.A4(n3120),
	.ZN(n3135));
   AOI22_X1 U3658 (.A1(REGISTERS[842]),
	.A2(n3570),
	.B1(REGISTERS[778]),
	.B2(n3569),
	.ZN(n3127));
   AOI22_X1 U3659 (.A1(REGISTERS[970]),
	.A2(FE_OFN46_n3572),
	.B1(REGISTERS[906]),
	.B2(FE_OFN6_n3571),
	.ZN(n3126));
   AOI22_X1 U3660 (.A1(REGISTERS[874]),
	.A2(FE_OFN4_n3574),
	.B1(REGISTERS[810]),
	.B2(FE_OFN133_n3573),
	.ZN(n3125));
   AOI22_X1 U3661 (.A1(REGISTERS[1002]),
	.A2(n3576),
	.B1(REGISTERS[938]),
	.B2(n3575),
	.ZN(n3124));
   NAND4_X1 U3662 (.A1(n3127),
	.A2(n3126),
	.A3(n3125),
	.A4(n3124),
	.ZN(n3133));
   AOI22_X1 U3663 (.A1(REGISTERS[586]),
	.A2(n3570),
	.B1(REGISTERS[522]),
	.B2(n3569),
	.ZN(n3131));
   AOI22_X1 U3664 (.A1(REGISTERS[714]),
	.A2(FE_OFN46_n3572),
	.B1(REGISTERS[650]),
	.B2(FE_OFN6_n3571),
	.ZN(n3130));
   AOI22_X1 U3665 (.A1(REGISTERS[618]),
	.A2(FE_OFN4_n3574),
	.B1(REGISTERS[554]),
	.B2(FE_OFN133_n3573),
	.ZN(n3129));
   AOI22_X1 U3666 (.A1(REGISTERS[746]),
	.A2(n3576),
	.B1(REGISTERS[682]),
	.B2(n3575),
	.ZN(n3128));
   NAND4_X1 U3667 (.A1(n3131),
	.A2(n3130),
	.A3(n3129),
	.A4(n3128),
	.ZN(n3132));
   AOI22_X1 U3668 (.A1(n3133),
	.A2(FE_OFN33_n3584),
	.B1(n3132),
	.B2(FE_OFN31_n3582),
	.ZN(n3134));
   OAI221_X1 U3669 (.A(n3134),
	.B1(FE_OFN38_n3588),
	.B2(n3136),
	.C1(n3586),
	.C2(n3135),
	.ZN(N117));
   AOI22_X1 U3670 (.A1(REGISTERS[331]),
	.A2(n3570),
	.B1(REGISTERS[267]),
	.B2(n3569),
	.ZN(n3140));
   AOI22_X1 U3671 (.A1(REGISTERS[459]),
	.A2(FE_OFN47_n3572),
	.B1(REGISTERS[395]),
	.B2(FE_OFN6_n3571),
	.ZN(n3139));
   AOI22_X1 U3672 (.A1(REGISTERS[363]),
	.A2(FE_OFN4_n3574),
	.B1(REGISTERS[299]),
	.B2(FE_OFN133_n3573),
	.ZN(n3138));
   AOI22_X1 U3673 (.A1(REGISTERS[491]),
	.A2(n3576),
	.B1(REGISTERS[427]),
	.B2(n3575),
	.ZN(n3137));
   AND4_X1 U3674 (.A1(n3140),
	.A2(n3139),
	.A3(n3138),
	.A4(n3137),
	.ZN(n3157));
   AOI22_X1 U3675 (.A1(REGISTERS[75]),
	.A2(n3570),
	.B1(REGISTERS[11]),
	.B2(n3569),
	.ZN(n3144));
   AOI22_X1 U3676 (.A1(REGISTERS[203]),
	.A2(FE_OFN47_n3572),
	.B1(REGISTERS[139]),
	.B2(FE_OFN6_n3571),
	.ZN(n3143));
   AOI22_X1 U3677 (.A1(REGISTERS[107]),
	.A2(FE_OFN4_n3574),
	.B1(REGISTERS[43]),
	.B2(FE_OFN133_n3573),
	.ZN(n3142));
   AOI22_X1 U3678 (.A1(REGISTERS[235]),
	.A2(n3576),
	.B1(REGISTERS[171]),
	.B2(n3575),
	.ZN(n3141));
   AND4_X1 U3679 (.A1(n3144),
	.A2(n3143),
	.A3(n3142),
	.A4(n3141),
	.ZN(n3156));
   AOI22_X1 U3680 (.A1(REGISTERS[843]),
	.A2(n3570),
	.B1(REGISTERS[779]),
	.B2(n3569),
	.ZN(n3148));
   AOI22_X1 U3681 (.A1(REGISTERS[971]),
	.A2(FE_OFN47_n3572),
	.B1(REGISTERS[907]),
	.B2(FE_OFN6_n3571),
	.ZN(n3147));
   AOI22_X1 U3682 (.A1(REGISTERS[875]),
	.A2(FE_OFN4_n3574),
	.B1(REGISTERS[811]),
	.B2(FE_OFN133_n3573),
	.ZN(n3146));
   AOI22_X1 U3683 (.A1(REGISTERS[1003]),
	.A2(n3576),
	.B1(REGISTERS[939]),
	.B2(n3575),
	.ZN(n3145));
   NAND4_X1 U3684 (.A1(n3148),
	.A2(n3147),
	.A3(n3146),
	.A4(n3145),
	.ZN(n3154));
   AOI22_X1 U3685 (.A1(REGISTERS[587]),
	.A2(n3570),
	.B1(REGISTERS[523]),
	.B2(n3569),
	.ZN(n3152));
   AOI22_X1 U3686 (.A1(REGISTERS[715]),
	.A2(FE_OFN47_n3572),
	.B1(REGISTERS[651]),
	.B2(FE_OFN6_n3571),
	.ZN(n3151));
   AOI22_X1 U3687 (.A1(REGISTERS[619]),
	.A2(FE_OFN4_n3574),
	.B1(REGISTERS[555]),
	.B2(FE_OFN133_n3573),
	.ZN(n3150));
   AOI22_X1 U3688 (.A1(REGISTERS[747]),
	.A2(n3576),
	.B1(REGISTERS[683]),
	.B2(n3575),
	.ZN(n3149));
   NAND4_X1 U3689 (.A1(n3152),
	.A2(n3151),
	.A3(n3150),
	.A4(n3149),
	.ZN(n3153));
   AOI22_X1 U3690 (.A1(n3154),
	.A2(FE_OFN33_n3584),
	.B1(n3153),
	.B2(FE_OFN31_n3582),
	.ZN(n3155));
   OAI221_X1 U3691 (.A(n3155),
	.B1(FE_OFN38_n3588),
	.B2(n3157),
	.C1(n3586),
	.C2(n3156),
	.ZN(N116));
   AOI22_X1 U3692 (.A1(REGISTERS[332]),
	.A2(n3570),
	.B1(REGISTERS[268]),
	.B2(FE_OFN108_n3569),
	.ZN(n3161));
   AOI22_X1 U3693 (.A1(REGISTERS[460]),
	.A2(n3572),
	.B1(REGISTERS[396]),
	.B2(n3571),
	.ZN(n3160));
   AOI22_X1 U3694 (.A1(REGISTERS[364]),
	.A2(n3574),
	.B1(REGISTERS[300]),
	.B2(n3573),
	.ZN(n3159));
   AOI22_X1 U3695 (.A1(REGISTERS[492]),
	.A2(n3576),
	.B1(REGISTERS[428]),
	.B2(n3575),
	.ZN(n3158));
   AND4_X1 U3696 (.A1(n3161),
	.A2(n3160),
	.A3(n3159),
	.A4(n3158),
	.ZN(n3178));
   AOI22_X1 U3697 (.A1(REGISTERS[76]),
	.A2(n3570),
	.B1(REGISTERS[12]),
	.B2(FE_OFN108_n3569),
	.ZN(n3165));
   AOI22_X1 U3698 (.A1(REGISTERS[204]),
	.A2(n3572),
	.B1(REGISTERS[140]),
	.B2(n3571),
	.ZN(n3164));
   AOI22_X1 U3699 (.A1(REGISTERS[108]),
	.A2(n3574),
	.B1(REGISTERS[44]),
	.B2(n3573),
	.ZN(n3163));
   AOI22_X1 U3700 (.A1(REGISTERS[236]),
	.A2(n3576),
	.B1(REGISTERS[172]),
	.B2(n3575),
	.ZN(n3162));
   AND4_X1 U3701 (.A1(n3165),
	.A2(n3164),
	.A3(n3163),
	.A4(n3162),
	.ZN(n3177));
   AOI22_X1 U3702 (.A1(REGISTERS[844]),
	.A2(n3570),
	.B1(REGISTERS[780]),
	.B2(n3569),
	.ZN(n3169));
   AOI22_X1 U3703 (.A1(REGISTERS[972]),
	.A2(FE_OFN46_n3572),
	.B1(REGISTERS[908]),
	.B2(FE_OFN6_n3571),
	.ZN(n3168));
   AOI22_X1 U3704 (.A1(REGISTERS[876]),
	.A2(FE_OFN4_n3574),
	.B1(REGISTERS[812]),
	.B2(FE_OFN133_n3573),
	.ZN(n3167));
   AOI22_X1 U3705 (.A1(REGISTERS[1004]),
	.A2(n3576),
	.B1(REGISTERS[940]),
	.B2(n3575),
	.ZN(n3166));
   NAND4_X1 U3706 (.A1(n3169),
	.A2(n3168),
	.A3(n3167),
	.A4(n3166),
	.ZN(n3175));
   AOI22_X1 U3707 (.A1(REGISTERS[588]),
	.A2(n3570),
	.B1(REGISTERS[524]),
	.B2(n3569),
	.ZN(n3173));
   AOI22_X1 U3708 (.A1(REGISTERS[716]),
	.A2(FE_OFN46_n3572),
	.B1(REGISTERS[652]),
	.B2(FE_OFN6_n3571),
	.ZN(n3172));
   AOI22_X1 U3709 (.A1(REGISTERS[620]),
	.A2(FE_OFN4_n3574),
	.B1(REGISTERS[556]),
	.B2(FE_OFN133_n3573),
	.ZN(n3171));
   AOI22_X1 U3710 (.A1(REGISTERS[748]),
	.A2(n3576),
	.B1(REGISTERS[684]),
	.B2(n3575),
	.ZN(n3170));
   NAND4_X1 U3711 (.A1(n3173),
	.A2(n3172),
	.A3(n3171),
	.A4(n3170),
	.ZN(n3174));
   AOI22_X1 U3712 (.A1(n3175),
	.A2(FE_OFN33_n3584),
	.B1(n3174),
	.B2(FE_OFN31_n3582),
	.ZN(n3176));
   OAI221_X1 U3713 (.A(n3176),
	.B1(FE_OFN38_n3588),
	.B2(n3178),
	.C1(n3586),
	.C2(n3177),
	.ZN(N115));
   AOI22_X1 U3714 (.A1(REGISTERS[333]),
	.A2(FE_OFN131_n3570),
	.B1(REGISTERS[269]),
	.B2(FE_OFN108_n3569),
	.ZN(n3182));
   AOI22_X1 U3715 (.A1(REGISTERS[461]),
	.A2(n3572),
	.B1(REGISTERS[397]),
	.B2(n3571),
	.ZN(n3181));
   AOI22_X1 U3716 (.A1(REGISTERS[365]),
	.A2(n3574),
	.B1(REGISTERS[301]),
	.B2(n3573),
	.ZN(n3180));
   AOI22_X1 U3717 (.A1(REGISTERS[493]),
	.A2(FE_OFN105_n3576),
	.B1(REGISTERS[429]),
	.B2(FE_OFN48_n3575),
	.ZN(n3179));
   AND4_X1 U3718 (.A1(n3182),
	.A2(n3181),
	.A3(n3180),
	.A4(n3179),
	.ZN(n3199));
   AOI22_X1 U3719 (.A1(REGISTERS[77]),
	.A2(FE_OFN131_n3570),
	.B1(REGISTERS[13]),
	.B2(FE_OFN108_n3569),
	.ZN(n3186));
   AOI22_X1 U3720 (.A1(REGISTERS[205]),
	.A2(n3572),
	.B1(REGISTERS[141]),
	.B2(n3571),
	.ZN(n3185));
   AOI22_X1 U3721 (.A1(REGISTERS[109]),
	.A2(n3574),
	.B1(REGISTERS[45]),
	.B2(n3573),
	.ZN(n3184));
   AOI22_X1 U3722 (.A1(REGISTERS[237]),
	.A2(FE_OFN105_n3576),
	.B1(REGISTERS[173]),
	.B2(FE_OFN48_n3575),
	.ZN(n3183));
   AND4_X1 U3723 (.A1(n3186),
	.A2(n3185),
	.A3(n3184),
	.A4(n3183),
	.ZN(n3198));
   AOI22_X1 U3724 (.A1(REGISTERS[845]),
	.A2(FE_OFN131_n3570),
	.B1(REGISTERS[781]),
	.B2(FE_OFN108_n3569),
	.ZN(n3190));
   AOI22_X1 U3725 (.A1(REGISTERS[973]),
	.A2(FE_OFN46_n3572),
	.B1(REGISTERS[909]),
	.B2(FE_OFN6_n3571),
	.ZN(n3189));
   AOI22_X1 U3726 (.A1(REGISTERS[877]),
	.A2(FE_OFN3_n3574),
	.B1(REGISTERS[813]),
	.B2(FE_OFN133_n3573),
	.ZN(n3188));
   AOI22_X1 U3727 (.A1(REGISTERS[1005]),
	.A2(FE_OFN105_n3576),
	.B1(REGISTERS[941]),
	.B2(FE_OFN48_n3575),
	.ZN(n3187));
   NAND4_X1 U3728 (.A1(n3190),
	.A2(n3189),
	.A3(n3188),
	.A4(n3187),
	.ZN(n3196));
   AOI22_X1 U3729 (.A1(REGISTERS[589]),
	.A2(FE_OFN131_n3570),
	.B1(REGISTERS[525]),
	.B2(FE_OFN108_n3569),
	.ZN(n3194));
   AOI22_X1 U3730 (.A1(REGISTERS[717]),
	.A2(FE_OFN46_n3572),
	.B1(REGISTERS[653]),
	.B2(FE_OFN6_n3571),
	.ZN(n3193));
   AOI22_X1 U3731 (.A1(REGISTERS[621]),
	.A2(FE_OFN3_n3574),
	.B1(REGISTERS[557]),
	.B2(FE_OFN133_n3573),
	.ZN(n3192));
   AOI22_X1 U3732 (.A1(REGISTERS[749]),
	.A2(FE_OFN105_n3576),
	.B1(REGISTERS[685]),
	.B2(FE_OFN48_n3575),
	.ZN(n3191));
   NAND4_X1 U3733 (.A1(n3194),
	.A2(n3193),
	.A3(n3192),
	.A4(n3191),
	.ZN(n3195));
   AOI22_X1 U3734 (.A1(n3196),
	.A2(FE_OFN33_n3584),
	.B1(n3195),
	.B2(FE_OFN31_n3582),
	.ZN(n3197));
   OAI221_X1 U3735 (.A(n3197),
	.B1(FE_OFN38_n3588),
	.B2(n3199),
	.C1(n3586),
	.C2(n3198),
	.ZN(N114));
   AOI22_X1 U3736 (.A1(REGISTERS[334]),
	.A2(FE_OFN132_n3570),
	.B1(REGISTERS[270]),
	.B2(FE_OFN109_n3569),
	.ZN(n3203));
   AOI22_X1 U3737 (.A1(REGISTERS[462]),
	.A2(FE_OFN47_n3572),
	.B1(REGISTERS[398]),
	.B2(FE_OFN6_n3571),
	.ZN(n3202));
   AOI22_X1 U3738 (.A1(REGISTERS[366]),
	.A2(FE_OFN4_n3574),
	.B1(REGISTERS[302]),
	.B2(FE_OFN133_n3573),
	.ZN(n3201));
   AOI22_X1 U3739 (.A1(REGISTERS[494]),
	.A2(FE_OFN107_n3576),
	.B1(REGISTERS[430]),
	.B2(FE_OFN50_n3575),
	.ZN(n3200));
   AND4_X1 U3740 (.A1(n3203),
	.A2(n3202),
	.A3(n3201),
	.A4(n3200),
	.ZN(n3220));
   AOI22_X1 U3741 (.A1(REGISTERS[78]),
	.A2(FE_OFN132_n3570),
	.B1(REGISTERS[14]),
	.B2(FE_OFN109_n3569),
	.ZN(n3207));
   AOI22_X1 U3742 (.A1(REGISTERS[206]),
	.A2(FE_OFN47_n3572),
	.B1(REGISTERS[142]),
	.B2(FE_OFN6_n3571),
	.ZN(n3206));
   AOI22_X1 U3743 (.A1(REGISTERS[110]),
	.A2(FE_OFN4_n3574),
	.B1(REGISTERS[46]),
	.B2(FE_OFN133_n3573),
	.ZN(n3205));
   AOI22_X1 U3744 (.A1(REGISTERS[238]),
	.A2(FE_OFN107_n3576),
	.B1(REGISTERS[174]),
	.B2(FE_OFN50_n3575),
	.ZN(n3204));
   AND4_X1 U3745 (.A1(n3207),
	.A2(n3206),
	.A3(n3205),
	.A4(n3204),
	.ZN(n3219));
   AOI22_X1 U3746 (.A1(REGISTERS[846]),
	.A2(FE_OFN132_n3570),
	.B1(REGISTERS[782]),
	.B2(FE_OFN109_n3569),
	.ZN(n3211));
   AOI22_X1 U3747 (.A1(REGISTERS[974]),
	.A2(FE_OFN47_n3572),
	.B1(REGISTERS[910]),
	.B2(FE_OFN7_n3571),
	.ZN(n3210));
   AOI22_X1 U3748 (.A1(REGISTERS[878]),
	.A2(FE_OFN5_n3574),
	.B1(REGISTERS[814]),
	.B2(FE_OFN134_n3573),
	.ZN(n3209));
   AOI22_X1 U3749 (.A1(REGISTERS[1006]),
	.A2(FE_OFN107_n3576),
	.B1(REGISTERS[942]),
	.B2(FE_OFN50_n3575),
	.ZN(n3208));
   NAND4_X1 U3750 (.A1(n3211),
	.A2(n3210),
	.A3(n3209),
	.A4(n3208),
	.ZN(n3217));
   AOI22_X1 U3751 (.A1(REGISTERS[590]),
	.A2(FE_OFN132_n3570),
	.B1(REGISTERS[526]),
	.B2(FE_OFN109_n3569),
	.ZN(n3215));
   AOI22_X1 U3752 (.A1(REGISTERS[718]),
	.A2(FE_OFN47_n3572),
	.B1(REGISTERS[654]),
	.B2(FE_OFN7_n3571),
	.ZN(n3214));
   AOI22_X1 U3753 (.A1(REGISTERS[622]),
	.A2(FE_OFN5_n3574),
	.B1(REGISTERS[558]),
	.B2(FE_OFN134_n3573),
	.ZN(n3213));
   AOI22_X1 U3754 (.A1(REGISTERS[750]),
	.A2(FE_OFN107_n3576),
	.B1(REGISTERS[686]),
	.B2(FE_OFN50_n3575),
	.ZN(n3212));
   NAND4_X1 U3755 (.A1(n3215),
	.A2(n3214),
	.A3(n3213),
	.A4(n3212),
	.ZN(n3216));
   AOI22_X1 U3756 (.A1(n3217),
	.A2(FE_OFN33_n3584),
	.B1(n3216),
	.B2(FE_OFN31_n3582),
	.ZN(n3218));
   OAI221_X1 U3757 (.A(n3218),
	.B1(FE_OFN38_n3588),
	.B2(n3220),
	.C1(n3586),
	.C2(n3219),
	.ZN(N113));
   AOI22_X1 U3758 (.A1(REGISTERS[335]),
	.A2(n3570),
	.B1(REGISTERS[271]),
	.B2(n3569),
	.ZN(n3224));
   AOI22_X1 U3759 (.A1(REGISTERS[463]),
	.A2(n3572),
	.B1(REGISTERS[399]),
	.B2(n3571),
	.ZN(n3223));
   AOI22_X1 U3760 (.A1(REGISTERS[367]),
	.A2(n3574),
	.B1(REGISTERS[303]),
	.B2(n3573),
	.ZN(n3222));
   AOI22_X1 U3761 (.A1(REGISTERS[495]),
	.A2(n3576),
	.B1(REGISTERS[431]),
	.B2(n3575),
	.ZN(n3221));
   AND4_X1 U3762 (.A1(n3224),
	.A2(n3223),
	.A3(n3222),
	.A4(n3221),
	.ZN(n3241));
   AOI22_X1 U3763 (.A1(REGISTERS[79]),
	.A2(n3570),
	.B1(REGISTERS[15]),
	.B2(FE_OFN108_n3569),
	.ZN(n3228));
   AOI22_X1 U3764 (.A1(REGISTERS[207]),
	.A2(n3572),
	.B1(REGISTERS[143]),
	.B2(n3571),
	.ZN(n3227));
   AOI22_X1 U3765 (.A1(REGISTERS[111]),
	.A2(n3574),
	.B1(REGISTERS[47]),
	.B2(n3573),
	.ZN(n3226));
   AOI22_X1 U3766 (.A1(REGISTERS[239]),
	.A2(n3576),
	.B1(REGISTERS[175]),
	.B2(n3575),
	.ZN(n3225));
   AND4_X1 U3767 (.A1(n3228),
	.A2(n3227),
	.A3(n3226),
	.A4(n3225),
	.ZN(n3240));
   AOI22_X1 U3768 (.A1(REGISTERS[847]),
	.A2(n3570),
	.B1(REGISTERS[783]),
	.B2(n3569),
	.ZN(n3232));
   AOI22_X1 U3769 (.A1(REGISTERS[975]),
	.A2(FE_OFN47_n3572),
	.B1(REGISTERS[911]),
	.B2(FE_OFN7_n3571),
	.ZN(n3231));
   AOI22_X1 U3770 (.A1(REGISTERS[879]),
	.A2(FE_OFN5_n3574),
	.B1(REGISTERS[815]),
	.B2(FE_OFN134_n3573),
	.ZN(n3230));
   AOI22_X1 U3771 (.A1(REGISTERS[1007]),
	.A2(FE_OFN107_n3576),
	.B1(REGISTERS[943]),
	.B2(FE_OFN50_n3575),
	.ZN(n3229));
   NAND4_X1 U3772 (.A1(n3232),
	.A2(n3231),
	.A3(n3230),
	.A4(n3229),
	.ZN(n3238));
   AOI22_X1 U3773 (.A1(REGISTERS[591]),
	.A2(n3570),
	.B1(REGISTERS[527]),
	.B2(n3569),
	.ZN(n3236));
   AOI22_X1 U3774 (.A1(REGISTERS[719]),
	.A2(FE_OFN47_n3572),
	.B1(REGISTERS[655]),
	.B2(FE_OFN7_n3571),
	.ZN(n3235));
   AOI22_X1 U3775 (.A1(REGISTERS[623]),
	.A2(FE_OFN5_n3574),
	.B1(REGISTERS[559]),
	.B2(FE_OFN134_n3573),
	.ZN(n3234));
   AOI22_X1 U3776 (.A1(REGISTERS[751]),
	.A2(FE_OFN107_n3576),
	.B1(REGISTERS[687]),
	.B2(FE_OFN50_n3575),
	.ZN(n3233));
   NAND4_X1 U3777 (.A1(n3236),
	.A2(n3235),
	.A3(n3234),
	.A4(n3233),
	.ZN(n3237));
   AOI22_X1 U3778 (.A1(n3238),
	.A2(FE_OFN33_n3584),
	.B1(n3237),
	.B2(FE_OFN31_n3582),
	.ZN(n3239));
   OAI221_X1 U3779 (.A(n3239),
	.B1(FE_OFN38_n3588),
	.B2(n3241),
	.C1(n3586),
	.C2(n3240),
	.ZN(N112));
   AOI22_X1 U3780 (.A1(REGISTERS[336]),
	.A2(n3570),
	.B1(REGISTERS[272]),
	.B2(n3569),
	.ZN(n3245));
   AOI22_X1 U3781 (.A1(REGISTERS[464]),
	.A2(FE_OFN47_n3572),
	.B1(REGISTERS[400]),
	.B2(FE_OFN6_n3571),
	.ZN(n3244));
   AOI22_X1 U3782 (.A1(REGISTERS[368]),
	.A2(FE_OFN4_n3574),
	.B1(REGISTERS[304]),
	.B2(FE_OFN133_n3573),
	.ZN(n3243));
   AOI22_X1 U3783 (.A1(REGISTERS[496]),
	.A2(n3576),
	.B1(REGISTERS[432]),
	.B2(n3575),
	.ZN(n3242));
   AND4_X1 U3784 (.A1(n3245),
	.A2(n3244),
	.A3(n3243),
	.A4(n3242),
	.ZN(n3262));
   AOI22_X1 U3785 (.A1(REGISTERS[80]),
	.A2(n3570),
	.B1(REGISTERS[16]),
	.B2(n3569),
	.ZN(n3249));
   AOI22_X1 U3786 (.A1(REGISTERS[208]),
	.A2(FE_OFN47_n3572),
	.B1(REGISTERS[144]),
	.B2(FE_OFN6_n3571),
	.ZN(n3248));
   AOI22_X1 U3787 (.A1(REGISTERS[112]),
	.A2(FE_OFN4_n3574),
	.B1(REGISTERS[48]),
	.B2(FE_OFN133_n3573),
	.ZN(n3247));
   AOI22_X1 U3788 (.A1(REGISTERS[240]),
	.A2(n3576),
	.B1(REGISTERS[176]),
	.B2(n3575),
	.ZN(n3246));
   AND4_X1 U3789 (.A1(n3249),
	.A2(n3248),
	.A3(n3247),
	.A4(n3246),
	.ZN(n3261));
   AOI22_X1 U3790 (.A1(REGISTERS[848]),
	.A2(n3570),
	.B1(REGISTERS[784]),
	.B2(n3569),
	.ZN(n3253));
   AOI22_X1 U3791 (.A1(REGISTERS[976]),
	.A2(FE_OFN47_n3572),
	.B1(REGISTERS[912]),
	.B2(FE_OFN7_n3571),
	.ZN(n3252));
   AOI22_X1 U3792 (.A1(REGISTERS[880]),
	.A2(FE_OFN4_n3574),
	.B1(REGISTERS[816]),
	.B2(FE_OFN133_n3573),
	.ZN(n3251));
   AOI22_X1 U3793 (.A1(REGISTERS[1008]),
	.A2(FE_OFN107_n3576),
	.B1(REGISTERS[944]),
	.B2(FE_OFN50_n3575),
	.ZN(n3250));
   NAND4_X1 U3794 (.A1(n3253),
	.A2(n3252),
	.A3(n3251),
	.A4(n3250),
	.ZN(n3259));
   AOI22_X1 U3795 (.A1(REGISTERS[592]),
	.A2(n3570),
	.B1(REGISTERS[528]),
	.B2(n3569),
	.ZN(n3257));
   AOI22_X1 U3796 (.A1(REGISTERS[720]),
	.A2(FE_OFN47_n3572),
	.B1(REGISTERS[656]),
	.B2(FE_OFN6_n3571),
	.ZN(n3256));
   AOI22_X1 U3797 (.A1(REGISTERS[624]),
	.A2(FE_OFN4_n3574),
	.B1(REGISTERS[560]),
	.B2(FE_OFN133_n3573),
	.ZN(n3255));
   AOI22_X1 U3798 (.A1(REGISTERS[752]),
	.A2(FE_OFN107_n3576),
	.B1(REGISTERS[688]),
	.B2(FE_OFN50_n3575),
	.ZN(n3254));
   NAND4_X1 U3799 (.A1(n3257),
	.A2(n3256),
	.A3(n3255),
	.A4(n3254),
	.ZN(n3258));
   AOI22_X1 U3800 (.A1(n3259),
	.A2(FE_OFN33_n3584),
	.B1(n3258),
	.B2(FE_OFN31_n3582),
	.ZN(n3260));
   OAI221_X1 U3801 (.A(n3260),
	.B1(FE_OFN38_n3588),
	.B2(n3262),
	.C1(n3586),
	.C2(n3261),
	.ZN(N111));
   AOI22_X1 U3802 (.A1(REGISTERS[337]),
	.A2(FE_OFN132_n3570),
	.B1(REGISTERS[273]),
	.B2(FE_OFN109_n3569),
	.ZN(n3266));
   AOI22_X1 U3803 (.A1(REGISTERS[465]),
	.A2(FE_OFN47_n3572),
	.B1(REGISTERS[401]),
	.B2(FE_OFN6_n3571),
	.ZN(n3265));
   AOI22_X1 U3804 (.A1(REGISTERS[369]),
	.A2(FE_OFN4_n3574),
	.B1(REGISTERS[305]),
	.B2(FE_OFN134_n3573),
	.ZN(n3264));
   AOI22_X1 U3805 (.A1(REGISTERS[497]),
	.A2(FE_OFN107_n3576),
	.B1(REGISTERS[433]),
	.B2(FE_OFN50_n3575),
	.ZN(n3263));
   AND4_X1 U3806 (.A1(n3266),
	.A2(n3265),
	.A3(n3264),
	.A4(n3263),
	.ZN(n3283));
   AOI22_X1 U3807 (.A1(REGISTERS[81]),
	.A2(FE_OFN132_n3570),
	.B1(REGISTERS[17]),
	.B2(FE_OFN109_n3569),
	.ZN(n3270));
   AOI22_X1 U3808 (.A1(REGISTERS[209]),
	.A2(FE_OFN47_n3572),
	.B1(REGISTERS[145]),
	.B2(FE_OFN7_n3571),
	.ZN(n3269));
   AOI22_X1 U3809 (.A1(REGISTERS[113]),
	.A2(FE_OFN4_n3574),
	.B1(REGISTERS[49]),
	.B2(FE_OFN134_n3573),
	.ZN(n3268));
   AOI22_X1 U3810 (.A1(REGISTERS[241]),
	.A2(FE_OFN107_n3576),
	.B1(REGISTERS[177]),
	.B2(FE_OFN50_n3575),
	.ZN(n3267));
   AND4_X1 U3811 (.A1(n3270),
	.A2(n3269),
	.A3(n3268),
	.A4(n3267),
	.ZN(n3282));
   AOI22_X1 U3812 (.A1(REGISTERS[849]),
	.A2(FE_OFN132_n3570),
	.B1(REGISTERS[785]),
	.B2(FE_OFN109_n3569),
	.ZN(n3274));
   AOI22_X1 U3813 (.A1(REGISTERS[977]),
	.A2(FE_OFN47_n3572),
	.B1(REGISTERS[913]),
	.B2(FE_OFN7_n3571),
	.ZN(n3273));
   AOI22_X1 U3814 (.A1(REGISTERS[881]),
	.A2(FE_OFN5_n3574),
	.B1(REGISTERS[817]),
	.B2(FE_OFN134_n3573),
	.ZN(n3272));
   AOI22_X1 U3815 (.A1(REGISTERS[1009]),
	.A2(FE_OFN107_n3576),
	.B1(REGISTERS[945]),
	.B2(FE_OFN49_n3575),
	.ZN(n3271));
   NAND4_X1 U3816 (.A1(n3274),
	.A2(n3273),
	.A3(n3272),
	.A4(n3271),
	.ZN(n3280));
   AOI22_X1 U3817 (.A1(REGISTERS[593]),
	.A2(FE_OFN132_n3570),
	.B1(REGISTERS[529]),
	.B2(FE_OFN109_n3569),
	.ZN(n3278));
   AOI22_X1 U3818 (.A1(REGISTERS[721]),
	.A2(FE_OFN47_n3572),
	.B1(REGISTERS[657]),
	.B2(FE_OFN7_n3571),
	.ZN(n3277));
   AOI22_X1 U3819 (.A1(REGISTERS[625]),
	.A2(FE_OFN5_n3574),
	.B1(REGISTERS[561]),
	.B2(FE_OFN134_n3573),
	.ZN(n3276));
   AOI22_X1 U3820 (.A1(REGISTERS[753]),
	.A2(FE_OFN107_n3576),
	.B1(REGISTERS[689]),
	.B2(FE_OFN49_n3575),
	.ZN(n3275));
   NAND4_X1 U3821 (.A1(n3278),
	.A2(n3277),
	.A3(n3276),
	.A4(n3275),
	.ZN(n3279));
   AOI22_X1 U3822 (.A1(n3280),
	.A2(FE_OFN33_n3584),
	.B1(n3279),
	.B2(FE_OFN31_n3582),
	.ZN(n3281));
   OAI221_X1 U3823 (.A(n3281),
	.B1(FE_OFN38_n3588),
	.B2(n3283),
	.C1(n3586),
	.C2(n3282),
	.ZN(N110));
   AOI22_X1 U3824 (.A1(REGISTERS[338]),
	.A2(FE_OFN131_n3570),
	.B1(REGISTERS[274]),
	.B2(FE_OFN108_n3569),
	.ZN(n3287));
   AOI22_X1 U3825 (.A1(REGISTERS[466]),
	.A2(n3572),
	.B1(REGISTERS[402]),
	.B2(n3571),
	.ZN(n3286));
   AOI22_X1 U3826 (.A1(REGISTERS[370]),
	.A2(n3574),
	.B1(REGISTERS[306]),
	.B2(n3573),
	.ZN(n3285));
   AOI22_X1 U3827 (.A1(REGISTERS[498]),
	.A2(FE_OFN105_n3576),
	.B1(REGISTERS[434]),
	.B2(FE_OFN48_n3575),
	.ZN(n3284));
   AND4_X1 U3828 (.A1(n3287),
	.A2(n3286),
	.A3(n3285),
	.A4(n3284),
	.ZN(n3304));
   AOI22_X1 U3829 (.A1(REGISTERS[82]),
	.A2(FE_OFN131_n3570),
	.B1(REGISTERS[18]),
	.B2(FE_OFN108_n3569),
	.ZN(n3291));
   AOI22_X1 U3830 (.A1(REGISTERS[210]),
	.A2(n3572),
	.B1(REGISTERS[146]),
	.B2(n3571),
	.ZN(n3290));
   AOI22_X1 U3831 (.A1(REGISTERS[114]),
	.A2(n3574),
	.B1(REGISTERS[50]),
	.B2(n3573),
	.ZN(n3289));
   AOI22_X1 U3832 (.A1(REGISTERS[242]),
	.A2(FE_OFN106_n3576),
	.B1(REGISTERS[178]),
	.B2(FE_OFN48_n3575),
	.ZN(n3288));
   AND4_X1 U3833 (.A1(n3291),
	.A2(n3290),
	.A3(n3289),
	.A4(n3288),
	.ZN(n3303));
   AOI22_X1 U3834 (.A1(REGISTERS[850]),
	.A2(FE_OFN131_n3570),
	.B1(REGISTERS[786]),
	.B2(FE_OFN108_n3569),
	.ZN(n3295));
   AOI22_X1 U3835 (.A1(REGISTERS[978]),
	.A2(FE_OFN46_n3572),
	.B1(REGISTERS[914]),
	.B2(n3571),
	.ZN(n3294));
   AOI22_X1 U3836 (.A1(REGISTERS[882]),
	.A2(n3574),
	.B1(REGISTERS[818]),
	.B2(n3573),
	.ZN(n3293));
   AOI22_X1 U3837 (.A1(REGISTERS[1010]),
	.A2(FE_OFN106_n3576),
	.B1(REGISTERS[946]),
	.B2(FE_OFN48_n3575),
	.ZN(n3292));
   NAND4_X1 U3838 (.A1(n3295),
	.A2(n3294),
	.A3(n3293),
	.A4(n3292),
	.ZN(n3301));
   AOI22_X1 U3839 (.A1(REGISTERS[594]),
	.A2(FE_OFN131_n3570),
	.B1(REGISTERS[530]),
	.B2(FE_OFN108_n3569),
	.ZN(n3299));
   AOI22_X1 U3840 (.A1(REGISTERS[722]),
	.A2(n3572),
	.B1(REGISTERS[658]),
	.B2(n3571),
	.ZN(n3298));
   AOI22_X1 U3841 (.A1(REGISTERS[626]),
	.A2(n3574),
	.B1(REGISTERS[562]),
	.B2(n3573),
	.ZN(n3297));
   AOI22_X1 U3842 (.A1(REGISTERS[754]),
	.A2(FE_OFN106_n3576),
	.B1(REGISTERS[690]),
	.B2(FE_OFN48_n3575),
	.ZN(n3296));
   NAND4_X1 U3843 (.A1(n3299),
	.A2(n3298),
	.A3(n3297),
	.A4(n3296),
	.ZN(n3300));
   AOI22_X1 U3844 (.A1(n3301),
	.A2(FE_OFN33_n3584),
	.B1(n3300),
	.B2(FE_OFN31_n3582),
	.ZN(n3302));
   OAI221_X1 U3845 (.A(n3302),
	.B1(FE_OFN38_n3588),
	.B2(n3304),
	.C1(n3586),
	.C2(n3303),
	.ZN(N109));
   AOI22_X1 U3846 (.A1(REGISTERS[339]),
	.A2(FE_OFN132_n3570),
	.B1(REGISTERS[275]),
	.B2(FE_OFN109_n3569),
	.ZN(n3308));
   AOI22_X1 U3847 (.A1(REGISTERS[467]),
	.A2(FE_OFN46_n3572),
	.B1(REGISTERS[403]),
	.B2(FE_OFN7_n3571),
	.ZN(n3307));
   AOI22_X1 U3848 (.A1(REGISTERS[371]),
	.A2(FE_OFN5_n3574),
	.B1(REGISTERS[307]),
	.B2(FE_OFN134_n3573),
	.ZN(n3306));
   AOI22_X1 U3849 (.A1(REGISTERS[499]),
	.A2(FE_OFN105_n3576),
	.B1(REGISTERS[435]),
	.B2(FE_OFN49_n3575),
	.ZN(n3305));
   AND4_X1 U3850 (.A1(n3308),
	.A2(n3307),
	.A3(n3306),
	.A4(n3305),
	.ZN(n3325));
   AOI22_X1 U3851 (.A1(REGISTERS[83]),
	.A2(FE_OFN132_n3570),
	.B1(REGISTERS[19]),
	.B2(FE_OFN109_n3569),
	.ZN(n3312));
   AOI22_X1 U3852 (.A1(REGISTERS[211]),
	.A2(FE_OFN46_n3572),
	.B1(REGISTERS[147]),
	.B2(FE_OFN7_n3571),
	.ZN(n3311));
   AOI22_X1 U3853 (.A1(REGISTERS[115]),
	.A2(FE_OFN5_n3574),
	.B1(REGISTERS[51]),
	.B2(FE_OFN134_n3573),
	.ZN(n3310));
   AOI22_X1 U3854 (.A1(REGISTERS[243]),
	.A2(FE_OFN105_n3576),
	.B1(REGISTERS[179]),
	.B2(FE_OFN49_n3575),
	.ZN(n3309));
   AND4_X1 U3855 (.A1(n3312),
	.A2(n3311),
	.A3(n3310),
	.A4(n3309),
	.ZN(n3324));
   AOI22_X1 U3856 (.A1(REGISTERS[851]),
	.A2(FE_OFN132_n3570),
	.B1(REGISTERS[787]),
	.B2(FE_OFN109_n3569),
	.ZN(n3316));
   AOI22_X1 U3857 (.A1(REGISTERS[979]),
	.A2(FE_OFN47_n3572),
	.B1(REGISTERS[915]),
	.B2(FE_OFN7_n3571),
	.ZN(n3315));
   AOI22_X1 U3858 (.A1(REGISTERS[883]),
	.A2(FE_OFN5_n3574),
	.B1(REGISTERS[819]),
	.B2(FE_OFN134_n3573),
	.ZN(n3314));
   AOI22_X1 U3859 (.A1(REGISTERS[1011]),
	.A2(FE_OFN107_n3576),
	.B1(REGISTERS[947]),
	.B2(FE_OFN49_n3575),
	.ZN(n3313));
   NAND4_X1 U3860 (.A1(n3316),
	.A2(n3315),
	.A3(n3314),
	.A4(n3313),
	.ZN(n3322));
   AOI22_X1 U3861 (.A1(REGISTERS[595]),
	.A2(FE_OFN132_n3570),
	.B1(REGISTERS[531]),
	.B2(FE_OFN109_n3569),
	.ZN(n3320));
   AOI22_X1 U3862 (.A1(REGISTERS[723]),
	.A2(FE_OFN47_n3572),
	.B1(REGISTERS[659]),
	.B2(FE_OFN7_n3571),
	.ZN(n3319));
   AOI22_X1 U3863 (.A1(REGISTERS[627]),
	.A2(FE_OFN5_n3574),
	.B1(REGISTERS[563]),
	.B2(FE_OFN134_n3573),
	.ZN(n3318));
   AOI22_X1 U3864 (.A1(REGISTERS[755]),
	.A2(FE_OFN107_n3576),
	.B1(REGISTERS[691]),
	.B2(FE_OFN49_n3575),
	.ZN(n3317));
   NAND4_X1 U3865 (.A1(n3320),
	.A2(n3319),
	.A3(n3318),
	.A4(n3317),
	.ZN(n3321));
   AOI22_X1 U3866 (.A1(n3322),
	.A2(FE_OFN33_n3584),
	.B1(n3321),
	.B2(FE_OFN31_n3582),
	.ZN(n3323));
   OAI221_X1 U3867 (.A(n3323),
	.B1(FE_OFN38_n3588),
	.B2(n3325),
	.C1(n3586),
	.C2(n3324),
	.ZN(N108));
   AOI22_X1 U3868 (.A1(REGISTERS[340]),
	.A2(FE_OFN131_n3570),
	.B1(REGISTERS[276]),
	.B2(FE_OFN108_n3569),
	.ZN(n3329));
   AOI22_X1 U3869 (.A1(REGISTERS[468]),
	.A2(n3572),
	.B1(REGISTERS[404]),
	.B2(n3571),
	.ZN(n3328));
   AOI22_X1 U3870 (.A1(REGISTERS[372]),
	.A2(n3574),
	.B1(REGISTERS[308]),
	.B2(n3573),
	.ZN(n3327));
   AOI22_X1 U3871 (.A1(REGISTERS[500]),
	.A2(FE_OFN106_n3576),
	.B1(REGISTERS[436]),
	.B2(FE_OFN48_n3575),
	.ZN(n3326));
   AND4_X1 U3872 (.A1(n3329),
	.A2(n3328),
	.A3(n3327),
	.A4(n3326),
	.ZN(n3346));
   AOI22_X1 U3873 (.A1(REGISTERS[84]),
	.A2(FE_OFN131_n3570),
	.B1(REGISTERS[20]),
	.B2(FE_OFN108_n3569),
	.ZN(n3333));
   AOI22_X1 U3874 (.A1(REGISTERS[212]),
	.A2(n3572),
	.B1(REGISTERS[148]),
	.B2(n3571),
	.ZN(n3332));
   AOI22_X1 U3875 (.A1(REGISTERS[116]),
	.A2(n3574),
	.B1(REGISTERS[52]),
	.B2(n3573),
	.ZN(n3331));
   AOI22_X1 U3876 (.A1(REGISTERS[244]),
	.A2(FE_OFN106_n3576),
	.B1(REGISTERS[180]),
	.B2(FE_OFN48_n3575),
	.ZN(n3330));
   AND4_X1 U3877 (.A1(n3333),
	.A2(n3332),
	.A3(n3331),
	.A4(n3330),
	.ZN(n3345));
   AOI22_X1 U3878 (.A1(REGISTERS[852]),
	.A2(FE_OFN131_n3570),
	.B1(REGISTERS[788]),
	.B2(FE_OFN108_n3569),
	.ZN(n3337));
   AOI22_X1 U3879 (.A1(REGISTERS[980]),
	.A2(FE_OFN46_n3572),
	.B1(REGISTERS[916]),
	.B2(n3571),
	.ZN(n3336));
   AOI22_X1 U3880 (.A1(REGISTERS[884]),
	.A2(n3574),
	.B1(REGISTERS[820]),
	.B2(n3573),
	.ZN(n3335));
   AOI22_X1 U3881 (.A1(REGISTERS[1012]),
	.A2(FE_OFN106_n3576),
	.B1(REGISTERS[948]),
	.B2(FE_OFN48_n3575),
	.ZN(n3334));
   NAND4_X1 U3882 (.A1(n3337),
	.A2(n3336),
	.A3(n3335),
	.A4(n3334),
	.ZN(n3343));
   AOI22_X1 U3883 (.A1(REGISTERS[596]),
	.A2(FE_OFN131_n3570),
	.B1(REGISTERS[532]),
	.B2(FE_OFN108_n3569),
	.ZN(n3341));
   AOI22_X1 U3884 (.A1(REGISTERS[724]),
	.A2(FE_OFN46_n3572),
	.B1(REGISTERS[660]),
	.B2(n3571),
	.ZN(n3340));
   AOI22_X1 U3885 (.A1(REGISTERS[628]),
	.A2(n3574),
	.B1(REGISTERS[564]),
	.B2(n3573),
	.ZN(n3339));
   AOI22_X1 U3886 (.A1(REGISTERS[756]),
	.A2(FE_OFN106_n3576),
	.B1(REGISTERS[692]),
	.B2(FE_OFN48_n3575),
	.ZN(n3338));
   NAND4_X1 U3887 (.A1(n3341),
	.A2(n3340),
	.A3(n3339),
	.A4(n3338),
	.ZN(n3342));
   AOI22_X1 U3888 (.A1(n3343),
	.A2(FE_OFN33_n3584),
	.B1(n3342),
	.B2(FE_OFN31_n3582),
	.ZN(n3344));
   OAI221_X1 U3889 (.A(n3344),
	.B1(FE_OFN38_n3588),
	.B2(n3346),
	.C1(n3586),
	.C2(n3345),
	.ZN(N107));
   AOI22_X1 U3890 (.A1(REGISTERS[341]),
	.A2(FE_OFN131_n3570),
	.B1(REGISTERS[277]),
	.B2(FE_OFN108_n3569),
	.ZN(n3350));
   AOI22_X1 U3891 (.A1(REGISTERS[469]),
	.A2(FE_OFN46_n3572),
	.B1(REGISTERS[405]),
	.B2(FE_OFN7_n3571),
	.ZN(n3349));
   AOI22_X1 U3892 (.A1(REGISTERS[373]),
	.A2(FE_OFN3_n3574),
	.B1(REGISTERS[309]),
	.B2(FE_OFN133_n3573),
	.ZN(n3348));
   AOI22_X1 U3893 (.A1(REGISTERS[501]),
	.A2(FE_OFN105_n3576),
	.B1(REGISTERS[437]),
	.B2(FE_OFN49_n3575),
	.ZN(n3347));
   AND4_X1 U3894 (.A1(n3350),
	.A2(n3349),
	.A3(n3348),
	.A4(n3347),
	.ZN(n3367));
   AOI22_X1 U3895 (.A1(REGISTERS[85]),
	.A2(FE_OFN132_n3570),
	.B1(REGISTERS[21]),
	.B2(FE_OFN109_n3569),
	.ZN(n3354));
   AOI22_X1 U3896 (.A1(REGISTERS[213]),
	.A2(FE_OFN46_n3572),
	.B1(REGISTERS[149]),
	.B2(FE_OFN7_n3571),
	.ZN(n3353));
   AOI22_X1 U3897 (.A1(REGISTERS[117]),
	.A2(FE_OFN5_n3574),
	.B1(REGISTERS[53]),
	.B2(FE_OFN134_n3573),
	.ZN(n3352));
   AOI22_X1 U3898 (.A1(REGISTERS[245]),
	.A2(FE_OFN105_n3576),
	.B1(REGISTERS[181]),
	.B2(FE_OFN49_n3575),
	.ZN(n3351));
   AND4_X1 U3899 (.A1(n3354),
	.A2(n3353),
	.A3(n3352),
	.A4(n3351),
	.ZN(n3366));
   AOI22_X1 U3900 (.A1(REGISTERS[853]),
	.A2(FE_OFN132_n3570),
	.B1(REGISTERS[789]),
	.B2(FE_OFN109_n3569),
	.ZN(n3358));
   AOI22_X1 U3901 (.A1(REGISTERS[981]),
	.A2(FE_OFN47_n3572),
	.B1(REGISTERS[917]),
	.B2(FE_OFN7_n3571),
	.ZN(n3357));
   AOI22_X1 U3902 (.A1(REGISTERS[885]),
	.A2(FE_OFN5_n3574),
	.B1(REGISTERS[821]),
	.B2(FE_OFN134_n3573),
	.ZN(n3356));
   AOI22_X1 U3903 (.A1(REGISTERS[1013]),
	.A2(FE_OFN105_n3576),
	.B1(REGISTERS[949]),
	.B2(FE_OFN49_n3575),
	.ZN(n3355));
   NAND4_X1 U3904 (.A1(n3358),
	.A2(n3357),
	.A3(n3356),
	.A4(n3355),
	.ZN(n3364));
   AOI22_X1 U3905 (.A1(REGISTERS[597]),
	.A2(FE_OFN132_n3570),
	.B1(REGISTERS[533]),
	.B2(FE_OFN109_n3569),
	.ZN(n3362));
   AOI22_X1 U3906 (.A1(REGISTERS[725]),
	.A2(FE_OFN47_n3572),
	.B1(REGISTERS[661]),
	.B2(FE_OFN7_n3571),
	.ZN(n3361));
   AOI22_X1 U3907 (.A1(REGISTERS[629]),
	.A2(FE_OFN5_n3574),
	.B1(REGISTERS[565]),
	.B2(FE_OFN134_n3573),
	.ZN(n3360));
   AOI22_X1 U3908 (.A1(REGISTERS[757]),
	.A2(FE_OFN105_n3576),
	.B1(REGISTERS[693]),
	.B2(FE_OFN49_n3575),
	.ZN(n3359));
   NAND4_X1 U3909 (.A1(n3362),
	.A2(n3361),
	.A3(n3360),
	.A4(n3359),
	.ZN(n3363));
   AOI22_X1 U3910 (.A1(n3364),
	.A2(FE_OFN33_n3584),
	.B1(n3363),
	.B2(FE_OFN31_n3582),
	.ZN(n3365));
   OAI221_X1 U3911 (.A(n3365),
	.B1(FE_OFN38_n3588),
	.B2(n3367),
	.C1(n3586),
	.C2(n3366),
	.ZN(N106));
   AOI22_X1 U3912 (.A1(REGISTERS[342]),
	.A2(FE_OFN131_n3570),
	.B1(REGISTERS[278]),
	.B2(FE_OFN108_n3569),
	.ZN(n3371));
   AOI22_X1 U3913 (.A1(REGISTERS[470]),
	.A2(FE_OFN46_n3572),
	.B1(REGISTERS[406]),
	.B2(FE_OFN7_n3571),
	.ZN(n3370));
   AOI22_X1 U3914 (.A1(REGISTERS[374]),
	.A2(FE_OFN3_n3574),
	.B1(REGISTERS[310]),
	.B2(FE_OFN133_n3573),
	.ZN(n3369));
   AOI22_X1 U3915 (.A1(REGISTERS[502]),
	.A2(FE_OFN105_n3576),
	.B1(REGISTERS[438]),
	.B2(FE_OFN49_n3575),
	.ZN(n3368));
   AND4_X1 U3916 (.A1(n3371),
	.A2(n3370),
	.A3(n3369),
	.A4(n3368),
	.ZN(n3388));
   AOI22_X1 U3917 (.A1(REGISTERS[86]),
	.A2(FE_OFN131_n3570),
	.B1(REGISTERS[22]),
	.B2(FE_OFN108_n3569),
	.ZN(n3375));
   AOI22_X1 U3918 (.A1(REGISTERS[214]),
	.A2(FE_OFN46_n3572),
	.B1(REGISTERS[150]),
	.B2(FE_OFN7_n3571),
	.ZN(n3374));
   AOI22_X1 U3919 (.A1(REGISTERS[118]),
	.A2(FE_OFN3_n3574),
	.B1(REGISTERS[54]),
	.B2(FE_OFN133_n3573),
	.ZN(n3373));
   AOI22_X1 U3920 (.A1(REGISTERS[246]),
	.A2(FE_OFN105_n3576),
	.B1(REGISTERS[182]),
	.B2(FE_OFN49_n3575),
	.ZN(n3372));
   AND4_X1 U3921 (.A1(n3375),
	.A2(n3374),
	.A3(n3373),
	.A4(n3372),
	.ZN(n3387));
   AOI22_X1 U3922 (.A1(REGISTERS[854]),
	.A2(FE_OFN132_n3570),
	.B1(REGISTERS[790]),
	.B2(FE_OFN109_n3569),
	.ZN(n3379));
   AOI22_X1 U3923 (.A1(REGISTERS[982]),
	.A2(FE_OFN47_n3572),
	.B1(REGISTERS[918]),
	.B2(FE_OFN7_n3571),
	.ZN(n3378));
   AOI22_X1 U3924 (.A1(REGISTERS[886]),
	.A2(FE_OFN5_n3574),
	.B1(REGISTERS[822]),
	.B2(FE_OFN134_n3573),
	.ZN(n3377));
   AOI22_X1 U3925 (.A1(REGISTERS[1014]),
	.A2(FE_OFN107_n3576),
	.B1(REGISTERS[950]),
	.B2(FE_OFN49_n3575),
	.ZN(n3376));
   NAND4_X1 U3926 (.A1(n3379),
	.A2(n3378),
	.A3(n3377),
	.A4(n3376),
	.ZN(n3385));
   AOI22_X1 U3927 (.A1(REGISTERS[598]),
	.A2(FE_OFN132_n3570),
	.B1(REGISTERS[534]),
	.B2(FE_OFN109_n3569),
	.ZN(n3383));
   AOI22_X1 U3928 (.A1(REGISTERS[726]),
	.A2(FE_OFN47_n3572),
	.B1(REGISTERS[662]),
	.B2(FE_OFN7_n3571),
	.ZN(n3382));
   AOI22_X1 U3929 (.A1(REGISTERS[630]),
	.A2(FE_OFN5_n3574),
	.B1(REGISTERS[566]),
	.B2(FE_OFN134_n3573),
	.ZN(n3381));
   AOI22_X1 U3930 (.A1(REGISTERS[758]),
	.A2(FE_OFN107_n3576),
	.B1(REGISTERS[694]),
	.B2(FE_OFN49_n3575),
	.ZN(n3380));
   NAND4_X1 U3931 (.A1(n3383),
	.A2(n3382),
	.A3(n3381),
	.A4(n3380),
	.ZN(n3384));
   AOI22_X1 U3932 (.A1(n3385),
	.A2(FE_OFN33_n3584),
	.B1(n3384),
	.B2(FE_OFN31_n3582),
	.ZN(n3386));
   OAI221_X1 U3933 (.A(n3386),
	.B1(FE_OFN38_n3588),
	.B2(n3388),
	.C1(n3586),
	.C2(n3387),
	.ZN(N105));
   AOI22_X1 U3934 (.A1(REGISTERS[343]),
	.A2(FE_OFN132_n3570),
	.B1(REGISTERS[279]),
	.B2(FE_OFN109_n3569),
	.ZN(n3392));
   AOI22_X1 U3935 (.A1(REGISTERS[471]),
	.A2(FE_OFN46_n3572),
	.B1(REGISTERS[407]),
	.B2(FE_OFN7_n3571),
	.ZN(n3391));
   AOI22_X1 U3936 (.A1(REGISTERS[375]),
	.A2(FE_OFN5_n3574),
	.B1(REGISTERS[311]),
	.B2(FE_OFN134_n3573),
	.ZN(n3390));
   AOI22_X1 U3937 (.A1(REGISTERS[503]),
	.A2(FE_OFN105_n3576),
	.B1(REGISTERS[439]),
	.B2(FE_OFN49_n3575),
	.ZN(n3389));
   AND4_X1 U3938 (.A1(n3392),
	.A2(n3391),
	.A3(n3390),
	.A4(n3389),
	.ZN(n3409));
   AOI22_X1 U3939 (.A1(REGISTERS[87]),
	.A2(FE_OFN132_n3570),
	.B1(REGISTERS[23]),
	.B2(FE_OFN109_n3569),
	.ZN(n3396));
   AOI22_X1 U3940 (.A1(REGISTERS[215]),
	.A2(FE_OFN46_n3572),
	.B1(REGISTERS[151]),
	.B2(FE_OFN7_n3571),
	.ZN(n3395));
   AOI22_X1 U3941 (.A1(REGISTERS[119]),
	.A2(FE_OFN5_n3574),
	.B1(REGISTERS[55]),
	.B2(FE_OFN134_n3573),
	.ZN(n3394));
   AOI22_X1 U3942 (.A1(REGISTERS[247]),
	.A2(FE_OFN105_n3576),
	.B1(REGISTERS[183]),
	.B2(FE_OFN49_n3575),
	.ZN(n3393));
   AND4_X1 U3943 (.A1(n3396),
	.A2(n3395),
	.A3(n3394),
	.A4(n3393),
	.ZN(n3408));
   AOI22_X1 U3944 (.A1(REGISTERS[855]),
	.A2(FE_OFN132_n3570),
	.B1(REGISTERS[791]),
	.B2(FE_OFN109_n3569),
	.ZN(n3400));
   AOI22_X1 U3945 (.A1(REGISTERS[983]),
	.A2(FE_OFN47_n3572),
	.B1(REGISTERS[919]),
	.B2(FE_OFN7_n3571),
	.ZN(n3399));
   AOI22_X1 U3946 (.A1(REGISTERS[887]),
	.A2(FE_OFN5_n3574),
	.B1(REGISTERS[823]),
	.B2(FE_OFN134_n3573),
	.ZN(n3398));
   AOI22_X1 U3947 (.A1(REGISTERS[1015]),
	.A2(FE_OFN107_n3576),
	.B1(REGISTERS[951]),
	.B2(FE_OFN49_n3575),
	.ZN(n3397));
   NAND4_X1 U3948 (.A1(n3400),
	.A2(n3399),
	.A3(n3398),
	.A4(n3397),
	.ZN(n3406));
   AOI22_X1 U3949 (.A1(REGISTERS[599]),
	.A2(FE_OFN132_n3570),
	.B1(REGISTERS[535]),
	.B2(FE_OFN109_n3569),
	.ZN(n3404));
   AOI22_X1 U3950 (.A1(REGISTERS[727]),
	.A2(FE_OFN47_n3572),
	.B1(REGISTERS[663]),
	.B2(FE_OFN7_n3571),
	.ZN(n3403));
   AOI22_X1 U3951 (.A1(REGISTERS[631]),
	.A2(FE_OFN5_n3574),
	.B1(REGISTERS[567]),
	.B2(FE_OFN134_n3573),
	.ZN(n3402));
   AOI22_X1 U3952 (.A1(REGISTERS[759]),
	.A2(FE_OFN107_n3576),
	.B1(REGISTERS[695]),
	.B2(FE_OFN49_n3575),
	.ZN(n3401));
   NAND4_X1 U3953 (.A1(n3404),
	.A2(n3403),
	.A3(n3402),
	.A4(n3401),
	.ZN(n3405));
   AOI22_X1 U3954 (.A1(n3406),
	.A2(FE_OFN33_n3584),
	.B1(n3405),
	.B2(FE_OFN31_n3582),
	.ZN(n3407));
   OAI221_X1 U3955 (.A(n3407),
	.B1(FE_OFN38_n3588),
	.B2(n3409),
	.C1(n3586),
	.C2(n3408),
	.ZN(N104));
   AOI22_X1 U3956 (.A1(REGISTERS[344]),
	.A2(FE_OFN131_n3570),
	.B1(REGISTERS[280]),
	.B2(FE_OFN108_n3569),
	.ZN(n3413));
   AOI22_X1 U3957 (.A1(REGISTERS[472]),
	.A2(n3572),
	.B1(REGISTERS[408]),
	.B2(n3571),
	.ZN(n3412));
   AOI22_X1 U3958 (.A1(REGISTERS[376]),
	.A2(n3574),
	.B1(REGISTERS[312]),
	.B2(n3573),
	.ZN(n3411));
   AOI22_X1 U3959 (.A1(REGISTERS[504]),
	.A2(FE_OFN106_n3576),
	.B1(REGISTERS[440]),
	.B2(FE_OFN48_n3575),
	.ZN(n3410));
   AND4_X1 U3960 (.A1(n3413),
	.A2(n3412),
	.A3(n3411),
	.A4(n3410),
	.ZN(n3430));
   AOI22_X1 U3961 (.A1(REGISTERS[88]),
	.A2(FE_OFN131_n3570),
	.B1(REGISTERS[24]),
	.B2(FE_OFN108_n3569),
	.ZN(n3417));
   AOI22_X1 U3962 (.A1(REGISTERS[216]),
	.A2(n3572),
	.B1(REGISTERS[152]),
	.B2(n3571),
	.ZN(n3416));
   AOI22_X1 U3963 (.A1(REGISTERS[120]),
	.A2(n3574),
	.B1(REGISTERS[56]),
	.B2(n3573),
	.ZN(n3415));
   AOI22_X1 U3964 (.A1(REGISTERS[248]),
	.A2(FE_OFN106_n3576),
	.B1(REGISTERS[184]),
	.B2(FE_OFN48_n3575),
	.ZN(n3414));
   AND4_X1 U3965 (.A1(n3417),
	.A2(n3416),
	.A3(n3415),
	.A4(n3414),
	.ZN(n3429));
   AOI22_X1 U3966 (.A1(REGISTERS[856]),
	.A2(FE_OFN131_n3570),
	.B1(REGISTERS[792]),
	.B2(FE_OFN108_n3569),
	.ZN(n3421));
   AOI22_X1 U3967 (.A1(REGISTERS[984]),
	.A2(FE_OFN46_n3572),
	.B1(REGISTERS[920]),
	.B2(n3571),
	.ZN(n3420));
   AOI22_X1 U3968 (.A1(REGISTERS[888]),
	.A2(n3574),
	.B1(REGISTERS[824]),
	.B2(n3573),
	.ZN(n3419));
   AOI22_X1 U3969 (.A1(REGISTERS[1016]),
	.A2(FE_OFN106_n3576),
	.B1(REGISTERS[952]),
	.B2(FE_OFN48_n3575),
	.ZN(n3418));
   NAND4_X1 U3970 (.A1(n3421),
	.A2(n3420),
	.A3(n3419),
	.A4(n3418),
	.ZN(n3427));
   AOI22_X1 U3971 (.A1(REGISTERS[600]),
	.A2(FE_OFN131_n3570),
	.B1(REGISTERS[536]),
	.B2(FE_OFN108_n3569),
	.ZN(n3425));
   AOI22_X1 U3972 (.A1(REGISTERS[728]),
	.A2(FE_OFN46_n3572),
	.B1(REGISTERS[664]),
	.B2(n3571),
	.ZN(n3424));
   AOI22_X1 U3973 (.A1(REGISTERS[632]),
	.A2(n3574),
	.B1(REGISTERS[568]),
	.B2(n3573),
	.ZN(n3423));
   AOI22_X1 U3974 (.A1(REGISTERS[760]),
	.A2(FE_OFN106_n3576),
	.B1(REGISTERS[696]),
	.B2(FE_OFN48_n3575),
	.ZN(n3422));
   NAND4_X1 U3975 (.A1(n3425),
	.A2(n3424),
	.A3(n3423),
	.A4(n3422),
	.ZN(n3426));
   AOI22_X1 U3976 (.A1(n3427),
	.A2(FE_OFN33_n3584),
	.B1(n3426),
	.B2(FE_OFN31_n3582),
	.ZN(n3428));
   OAI221_X1 U3977 (.A(n3428),
	.B1(FE_OFN38_n3588),
	.B2(n3430),
	.C1(n3586),
	.C2(n3429),
	.ZN(N103));
   AOI22_X1 U3978 (.A1(REGISTERS[345]),
	.A2(FE_OFN132_n3570),
	.B1(REGISTERS[281]),
	.B2(FE_OFN109_n3569),
	.ZN(n3434));
   AOI22_X1 U3979 (.A1(REGISTERS[473]),
	.A2(FE_OFN46_n3572),
	.B1(REGISTERS[409]),
	.B2(FE_OFN7_n3571),
	.ZN(n3433));
   AOI22_X1 U3980 (.A1(REGISTERS[377]),
	.A2(FE_OFN5_n3574),
	.B1(REGISTERS[313]),
	.B2(FE_OFN134_n3573),
	.ZN(n3432));
   AOI22_X1 U3981 (.A1(REGISTERS[505]),
	.A2(FE_OFN105_n3576),
	.B1(REGISTERS[441]),
	.B2(FE_OFN49_n3575),
	.ZN(n3431));
   AND4_X1 U3982 (.A1(n3434),
	.A2(n3433),
	.A3(n3432),
	.A4(n3431),
	.ZN(n3451));
   AOI22_X1 U3983 (.A1(REGISTERS[89]),
	.A2(FE_OFN132_n3570),
	.B1(REGISTERS[25]),
	.B2(FE_OFN109_n3569),
	.ZN(n3438));
   AOI22_X1 U3984 (.A1(REGISTERS[217]),
	.A2(FE_OFN46_n3572),
	.B1(REGISTERS[153]),
	.B2(FE_OFN7_n3571),
	.ZN(n3437));
   AOI22_X1 U3985 (.A1(REGISTERS[121]),
	.A2(FE_OFN5_n3574),
	.B1(REGISTERS[57]),
	.B2(FE_OFN134_n3573),
	.ZN(n3436));
   AOI22_X1 U3986 (.A1(REGISTERS[249]),
	.A2(FE_OFN105_n3576),
	.B1(REGISTERS[185]),
	.B2(FE_OFN49_n3575),
	.ZN(n3435));
   AND4_X1 U3987 (.A1(n3438),
	.A2(n3437),
	.A3(n3436),
	.A4(n3435),
	.ZN(n3450));
   AOI22_X1 U3988 (.A1(REGISTERS[857]),
	.A2(FE_OFN132_n3570),
	.B1(REGISTERS[793]),
	.B2(FE_OFN109_n3569),
	.ZN(n3442));
   AOI22_X1 U3989 (.A1(REGISTERS[985]),
	.A2(FE_OFN47_n3572),
	.B1(REGISTERS[921]),
	.B2(FE_OFN7_n3571),
	.ZN(n3441));
   AOI22_X1 U3990 (.A1(REGISTERS[889]),
	.A2(FE_OFN5_n3574),
	.B1(REGISTERS[825]),
	.B2(FE_OFN134_n3573),
	.ZN(n3440));
   AOI22_X1 U3991 (.A1(REGISTERS[1017]),
	.A2(FE_OFN107_n3576),
	.B1(REGISTERS[953]),
	.B2(FE_OFN49_n3575),
	.ZN(n3439));
   NAND4_X1 U3992 (.A1(n3442),
	.A2(n3441),
	.A3(n3440),
	.A4(n3439),
	.ZN(n3448));
   AOI22_X1 U3993 (.A1(REGISTERS[601]),
	.A2(FE_OFN132_n3570),
	.B1(REGISTERS[537]),
	.B2(FE_OFN109_n3569),
	.ZN(n3446));
   AOI22_X1 U3994 (.A1(REGISTERS[729]),
	.A2(FE_OFN47_n3572),
	.B1(REGISTERS[665]),
	.B2(FE_OFN7_n3571),
	.ZN(n3445));
   AOI22_X1 U3995 (.A1(REGISTERS[633]),
	.A2(FE_OFN5_n3574),
	.B1(REGISTERS[569]),
	.B2(FE_OFN134_n3573),
	.ZN(n3444));
   AOI22_X1 U3996 (.A1(REGISTERS[761]),
	.A2(FE_OFN107_n3576),
	.B1(REGISTERS[697]),
	.B2(FE_OFN49_n3575),
	.ZN(n3443));
   NAND4_X1 U3997 (.A1(n3446),
	.A2(n3445),
	.A3(n3444),
	.A4(n3443),
	.ZN(n3447));
   AOI22_X1 U3998 (.A1(n3448),
	.A2(FE_OFN33_n3584),
	.B1(n3447),
	.B2(FE_OFN31_n3582),
	.ZN(n3449));
   OAI221_X1 U3999 (.A(n3449),
	.B1(FE_OFN38_n3588),
	.B2(n3451),
	.C1(n3586),
	.C2(n3450),
	.ZN(N102));
   AOI22_X1 U4000 (.A1(REGISTERS[346]),
	.A2(FE_OFN131_n3570),
	.B1(REGISTERS[282]),
	.B2(FE_OFN108_n3569),
	.ZN(n3455));
   AOI22_X1 U4001 (.A1(REGISTERS[474]),
	.A2(n3572),
	.B1(REGISTERS[410]),
	.B2(n3571),
	.ZN(n3454));
   AOI22_X1 U4002 (.A1(REGISTERS[378]),
	.A2(n3574),
	.B1(REGISTERS[314]),
	.B2(n3573),
	.ZN(n3453));
   AOI22_X1 U4003 (.A1(REGISTERS[506]),
	.A2(FE_OFN106_n3576),
	.B1(REGISTERS[442]),
	.B2(FE_OFN48_n3575),
	.ZN(n3452));
   AND4_X1 U4004 (.A1(n3455),
	.A2(n3454),
	.A3(n3453),
	.A4(n3452),
	.ZN(n3472));
   AOI22_X1 U4005 (.A1(REGISTERS[90]),
	.A2(FE_OFN131_n3570),
	.B1(REGISTERS[26]),
	.B2(FE_OFN108_n3569),
	.ZN(n3459));
   AOI22_X1 U4006 (.A1(REGISTERS[218]),
	.A2(n3572),
	.B1(REGISTERS[154]),
	.B2(n3571),
	.ZN(n3458));
   AOI22_X1 U4007 (.A1(REGISTERS[122]),
	.A2(n3574),
	.B1(REGISTERS[58]),
	.B2(n3573),
	.ZN(n3457));
   AOI22_X1 U4008 (.A1(REGISTERS[250]),
	.A2(FE_OFN106_n3576),
	.B1(REGISTERS[186]),
	.B2(FE_OFN48_n3575),
	.ZN(n3456));
   AND4_X1 U4009 (.A1(n3459),
	.A2(n3458),
	.A3(n3457),
	.A4(n3456),
	.ZN(n3471));
   AOI22_X1 U4010 (.A1(REGISTERS[858]),
	.A2(FE_OFN131_n3570),
	.B1(REGISTERS[794]),
	.B2(FE_OFN108_n3569),
	.ZN(n3463));
   AOI22_X1 U4011 (.A1(REGISTERS[986]),
	.A2(FE_OFN46_n3572),
	.B1(REGISTERS[922]),
	.B2(n3571),
	.ZN(n3462));
   AOI22_X1 U4012 (.A1(REGISTERS[890]),
	.A2(n3574),
	.B1(REGISTERS[826]),
	.B2(n3573),
	.ZN(n3461));
   AOI22_X1 U4013 (.A1(REGISTERS[1018]),
	.A2(FE_OFN106_n3576),
	.B1(REGISTERS[954]),
	.B2(FE_OFN48_n3575),
	.ZN(n3460));
   NAND4_X1 U4014 (.A1(n3463),
	.A2(n3462),
	.A3(n3461),
	.A4(n3460),
	.ZN(n3469));
   AOI22_X1 U4015 (.A1(REGISTERS[602]),
	.A2(FE_OFN131_n3570),
	.B1(REGISTERS[538]),
	.B2(FE_OFN108_n3569),
	.ZN(n3467));
   AOI22_X1 U4016 (.A1(REGISTERS[730]),
	.A2(FE_OFN46_n3572),
	.B1(REGISTERS[666]),
	.B2(n3571),
	.ZN(n3466));
   AOI22_X1 U4017 (.A1(REGISTERS[634]),
	.A2(n3574),
	.B1(REGISTERS[570]),
	.B2(n3573),
	.ZN(n3465));
   AOI22_X1 U4018 (.A1(REGISTERS[762]),
	.A2(FE_OFN106_n3576),
	.B1(REGISTERS[698]),
	.B2(FE_OFN48_n3575),
	.ZN(n3464));
   NAND4_X1 U4019 (.A1(n3467),
	.A2(n3466),
	.A3(n3465),
	.A4(n3464),
	.ZN(n3468));
   AOI22_X1 U4020 (.A1(n3469),
	.A2(FE_OFN33_n3584),
	.B1(n3468),
	.B2(FE_OFN31_n3582),
	.ZN(n3470));
   OAI221_X1 U4021 (.A(n3470),
	.B1(FE_OFN38_n3588),
	.B2(n3472),
	.C1(n3586),
	.C2(n3471),
	.ZN(N101));
   AOI22_X1 U4022 (.A1(REGISTERS[347]),
	.A2(FE_OFN132_n3570),
	.B1(REGISTERS[283]),
	.B2(FE_OFN109_n3569),
	.ZN(n3476));
   AOI22_X1 U4023 (.A1(REGISTERS[475]),
	.A2(FE_OFN47_n3572),
	.B1(REGISTERS[411]),
	.B2(FE_OFN7_n3571),
	.ZN(n3475));
   AOI22_X1 U4024 (.A1(REGISTERS[379]),
	.A2(FE_OFN4_n3574),
	.B1(REGISTERS[315]),
	.B2(FE_OFN134_n3573),
	.ZN(n3474));
   AOI22_X1 U4025 (.A1(REGISTERS[507]),
	.A2(FE_OFN107_n3576),
	.B1(REGISTERS[443]),
	.B2(FE_OFN50_n3575),
	.ZN(n3473));
   AND4_X1 U4026 (.A1(n3476),
	.A2(n3475),
	.A3(n3474),
	.A4(n3473),
	.ZN(n3493));
   AOI22_X1 U4027 (.A1(REGISTERS[91]),
	.A2(FE_OFN132_n3570),
	.B1(REGISTERS[27]),
	.B2(FE_OFN109_n3569),
	.ZN(n3480));
   AOI22_X1 U4028 (.A1(REGISTERS[219]),
	.A2(FE_OFN47_n3572),
	.B1(REGISTERS[155]),
	.B2(FE_OFN7_n3571),
	.ZN(n3479));
   AOI22_X1 U4029 (.A1(REGISTERS[123]),
	.A2(FE_OFN4_n3574),
	.B1(REGISTERS[59]),
	.B2(FE_OFN134_n3573),
	.ZN(n3478));
   AOI22_X1 U4030 (.A1(REGISTERS[251]),
	.A2(FE_OFN107_n3576),
	.B1(REGISTERS[187]),
	.B2(FE_OFN50_n3575),
	.ZN(n3477));
   AND4_X1 U4031 (.A1(n3480),
	.A2(n3479),
	.A3(n3478),
	.A4(n3477),
	.ZN(n3492));
   AOI22_X1 U4032 (.A1(REGISTERS[859]),
	.A2(FE_OFN132_n3570),
	.B1(REGISTERS[795]),
	.B2(FE_OFN109_n3569),
	.ZN(n3484));
   AOI22_X1 U4033 (.A1(REGISTERS[987]),
	.A2(FE_OFN47_n3572),
	.B1(REGISTERS[923]),
	.B2(FE_OFN7_n3571),
	.ZN(n3483));
   AOI22_X1 U4034 (.A1(REGISTERS[891]),
	.A2(FE_OFN5_n3574),
	.B1(REGISTERS[827]),
	.B2(FE_OFN134_n3573),
	.ZN(n3482));
   AOI22_X1 U4035 (.A1(REGISTERS[1019]),
	.A2(FE_OFN107_n3576),
	.B1(REGISTERS[955]),
	.B2(FE_OFN49_n3575),
	.ZN(n3481));
   NAND4_X1 U4036 (.A1(n3484),
	.A2(n3483),
	.A3(n3482),
	.A4(n3481),
	.ZN(n3490));
   AOI22_X1 U4037 (.A1(REGISTERS[603]),
	.A2(FE_OFN132_n3570),
	.B1(REGISTERS[539]),
	.B2(FE_OFN109_n3569),
	.ZN(n3488));
   AOI22_X1 U4038 (.A1(REGISTERS[731]),
	.A2(FE_OFN47_n3572),
	.B1(REGISTERS[667]),
	.B2(FE_OFN7_n3571),
	.ZN(n3487));
   AOI22_X1 U4039 (.A1(REGISTERS[635]),
	.A2(FE_OFN5_n3574),
	.B1(REGISTERS[571]),
	.B2(FE_OFN134_n3573),
	.ZN(n3486));
   AOI22_X1 U4040 (.A1(REGISTERS[763]),
	.A2(FE_OFN107_n3576),
	.B1(REGISTERS[699]),
	.B2(FE_OFN49_n3575),
	.ZN(n3485));
   NAND4_X1 U4041 (.A1(n3488),
	.A2(n3487),
	.A3(n3486),
	.A4(n3485),
	.ZN(n3489));
   AOI22_X1 U4042 (.A1(n3490),
	.A2(FE_OFN33_n3584),
	.B1(n3489),
	.B2(FE_OFN31_n3582),
	.ZN(n3491));
   OAI221_X1 U4043 (.A(n3491),
	.B1(FE_OFN38_n3588),
	.B2(n3493),
	.C1(n3586),
	.C2(n3492),
	.ZN(N100));
   AOI22_X1 U4044 (.A1(REGISTERS[348]),
	.A2(FE_OFN131_n3570),
	.B1(REGISTERS[284]),
	.B2(FE_OFN108_n3569),
	.ZN(n3497));
   AOI22_X1 U4045 (.A1(REGISTERS[476]),
	.A2(FE_OFN46_n3572),
	.B1(REGISTERS[412]),
	.B2(FE_OFN7_n3571),
	.ZN(n3496));
   AOI22_X1 U4046 (.A1(REGISTERS[380]),
	.A2(FE_OFN3_n3574),
	.B1(REGISTERS[316]),
	.B2(FE_OFN133_n3573),
	.ZN(n3495));
   AOI22_X1 U4047 (.A1(REGISTERS[508]),
	.A2(FE_OFN105_n3576),
	.B1(REGISTERS[444]),
	.B2(FE_OFN49_n3575),
	.ZN(n3494));
   AND4_X1 U4048 (.A1(n3497),
	.A2(n3496),
	.A3(n3495),
	.A4(n3494),
	.ZN(n3514));
   AOI22_X1 U4049 (.A1(REGISTERS[92]),
	.A2(FE_OFN131_n3570),
	.B1(REGISTERS[28]),
	.B2(FE_OFN108_n3569),
	.ZN(n3501));
   AOI22_X1 U4050 (.A1(REGISTERS[220]),
	.A2(FE_OFN46_n3572),
	.B1(REGISTERS[156]),
	.B2(FE_OFN7_n3571),
	.ZN(n3500));
   AOI22_X1 U4051 (.A1(REGISTERS[124]),
	.A2(FE_OFN3_n3574),
	.B1(REGISTERS[60]),
	.B2(FE_OFN133_n3573),
	.ZN(n3499));
   AOI22_X1 U4052 (.A1(REGISTERS[252]),
	.A2(FE_OFN105_n3576),
	.B1(REGISTERS[188]),
	.B2(FE_OFN49_n3575),
	.ZN(n3498));
   AND4_X1 U4053 (.A1(n3501),
	.A2(n3500),
	.A3(n3499),
	.A4(n3498),
	.ZN(n3513));
   AOI22_X1 U4054 (.A1(REGISTERS[860]),
	.A2(FE_OFN132_n3570),
	.B1(REGISTERS[796]),
	.B2(FE_OFN109_n3569),
	.ZN(n3505));
   AOI22_X1 U4055 (.A1(REGISTERS[988]),
	.A2(FE_OFN47_n3572),
	.B1(REGISTERS[924]),
	.B2(FE_OFN7_n3571),
	.ZN(n3504));
   AOI22_X1 U4056 (.A1(REGISTERS[892]),
	.A2(FE_OFN5_n3574),
	.B1(REGISTERS[828]),
	.B2(FE_OFN134_n3573),
	.ZN(n3503));
   AOI22_X1 U4057 (.A1(REGISTERS[1020]),
	.A2(FE_OFN107_n3576),
	.B1(REGISTERS[956]),
	.B2(FE_OFN49_n3575),
	.ZN(n3502));
   NAND4_X1 U4058 (.A1(n3505),
	.A2(n3504),
	.A3(n3503),
	.A4(n3502),
	.ZN(n3511));
   AOI22_X1 U4059 (.A1(REGISTERS[604]),
	.A2(FE_OFN132_n3570),
	.B1(REGISTERS[540]),
	.B2(FE_OFN109_n3569),
	.ZN(n3509));
   AOI22_X1 U4060 (.A1(REGISTERS[732]),
	.A2(FE_OFN47_n3572),
	.B1(REGISTERS[668]),
	.B2(FE_OFN7_n3571),
	.ZN(n3508));
   AOI22_X1 U4061 (.A1(REGISTERS[636]),
	.A2(FE_OFN5_n3574),
	.B1(REGISTERS[572]),
	.B2(FE_OFN134_n3573),
	.ZN(n3507));
   AOI22_X1 U4062 (.A1(REGISTERS[764]),
	.A2(FE_OFN107_n3576),
	.B1(REGISTERS[700]),
	.B2(FE_OFN49_n3575),
	.ZN(n3506));
   NAND4_X1 U4063 (.A1(n3509),
	.A2(n3508),
	.A3(n3507),
	.A4(n3506),
	.ZN(n3510));
   AOI22_X1 U4064 (.A1(n3511),
	.A2(FE_OFN33_n3584),
	.B1(n3510),
	.B2(FE_OFN31_n3582),
	.ZN(n3512));
   OAI221_X1 U4065 (.A(n3512),
	.B1(FE_OFN38_n3588),
	.B2(n3514),
	.C1(n3586),
	.C2(n3513),
	.ZN(N99));
   AOI22_X1 U4066 (.A1(REGISTERS[349]),
	.A2(FE_OFN131_n3570),
	.B1(REGISTERS[285]),
	.B2(FE_OFN108_n3569),
	.ZN(n3518));
   AOI22_X1 U4067 (.A1(REGISTERS[477]),
	.A2(FE_OFN46_n3572),
	.B1(REGISTERS[413]),
	.B2(FE_OFN6_n3571),
	.ZN(n3517));
   AOI22_X1 U4068 (.A1(REGISTERS[381]),
	.A2(FE_OFN3_n3574),
	.B1(REGISTERS[317]),
	.B2(FE_OFN133_n3573),
	.ZN(n3516));
   AOI22_X1 U4069 (.A1(REGISTERS[509]),
	.A2(FE_OFN105_n3576),
	.B1(REGISTERS[445]),
	.B2(FE_OFN48_n3575),
	.ZN(n3515));
   AND4_X1 U4070 (.A1(n3518),
	.A2(n3517),
	.A3(n3516),
	.A4(n3515),
	.ZN(n3535));
   AOI22_X1 U4071 (.A1(REGISTERS[93]),
	.A2(FE_OFN131_n3570),
	.B1(REGISTERS[29]),
	.B2(FE_OFN108_n3569),
	.ZN(n3522));
   AOI22_X1 U4072 (.A1(REGISTERS[221]),
	.A2(FE_OFN46_n3572),
	.B1(REGISTERS[157]),
	.B2(FE_OFN6_n3571),
	.ZN(n3521));
   AOI22_X1 U4073 (.A1(REGISTERS[125]),
	.A2(FE_OFN3_n3574),
	.B1(REGISTERS[61]),
	.B2(FE_OFN133_n3573),
	.ZN(n3520));
   AOI22_X1 U4074 (.A1(REGISTERS[253]),
	.A2(FE_OFN105_n3576),
	.B1(REGISTERS[189]),
	.B2(FE_OFN48_n3575),
	.ZN(n3519));
   AND4_X1 U4075 (.A1(n3522),
	.A2(n3521),
	.A3(n3520),
	.A4(n3519),
	.ZN(n3534));
   AOI22_X1 U4076 (.A1(REGISTERS[861]),
	.A2(FE_OFN131_n3570),
	.B1(REGISTERS[797]),
	.B2(FE_OFN108_n3569),
	.ZN(n3526));
   AOI22_X1 U4077 (.A1(REGISTERS[989]),
	.A2(FE_OFN46_n3572),
	.B1(REGISTERS[925]),
	.B2(FE_OFN6_n3571),
	.ZN(n3525));
   AOI22_X1 U4078 (.A1(REGISTERS[893]),
	.A2(FE_OFN3_n3574),
	.B1(REGISTERS[829]),
	.B2(FE_OFN133_n3573),
	.ZN(n3524));
   AOI22_X1 U4079 (.A1(REGISTERS[1021]),
	.A2(FE_OFN105_n3576),
	.B1(REGISTERS[957]),
	.B2(FE_OFN49_n3575),
	.ZN(n3523));
   NAND4_X1 U4080 (.A1(n3526),
	.A2(n3525),
	.A3(n3524),
	.A4(n3523),
	.ZN(n3532));
   AOI22_X1 U4081 (.A1(REGISTERS[605]),
	.A2(FE_OFN131_n3570),
	.B1(REGISTERS[541]),
	.B2(FE_OFN108_n3569),
	.ZN(n3530));
   AOI22_X1 U4082 (.A1(REGISTERS[733]),
	.A2(FE_OFN46_n3572),
	.B1(REGISTERS[669]),
	.B2(FE_OFN6_n3571),
	.ZN(n3529));
   AOI22_X1 U4083 (.A1(REGISTERS[637]),
	.A2(FE_OFN3_n3574),
	.B1(REGISTERS[573]),
	.B2(FE_OFN133_n3573),
	.ZN(n3528));
   AOI22_X1 U4084 (.A1(REGISTERS[765]),
	.A2(FE_OFN105_n3576),
	.B1(REGISTERS[701]),
	.B2(FE_OFN48_n3575),
	.ZN(n3527));
   NAND4_X1 U4085 (.A1(n3530),
	.A2(n3529),
	.A3(n3528),
	.A4(n3527),
	.ZN(n3531));
   AOI22_X1 U4086 (.A1(n3532),
	.A2(FE_OFN33_n3584),
	.B1(n3531),
	.B2(FE_OFN31_n3582),
	.ZN(n3533));
   OAI221_X1 U4087 (.A(n3533),
	.B1(FE_OFN38_n3588),
	.B2(n3535),
	.C1(n3586),
	.C2(n3534),
	.ZN(N98));
   AOI22_X1 U4088 (.A1(REGISTERS[350]),
	.A2(FE_OFN131_n3570),
	.B1(REGISTERS[286]),
	.B2(FE_OFN108_n3569),
	.ZN(n3539));
   AOI22_X1 U4089 (.A1(REGISTERS[478]),
	.A2(FE_OFN46_n3572),
	.B1(REGISTERS[414]),
	.B2(FE_OFN7_n3571),
	.ZN(n3538));
   AOI22_X1 U4090 (.A1(REGISTERS[382]),
	.A2(FE_OFN3_n3574),
	.B1(REGISTERS[318]),
	.B2(FE_OFN133_n3573),
	.ZN(n3537));
   AOI22_X1 U4091 (.A1(REGISTERS[510]),
	.A2(FE_OFN105_n3576),
	.B1(REGISTERS[446]),
	.B2(FE_OFN49_n3575),
	.ZN(n3536));
   AND4_X1 U4092 (.A1(n3539),
	.A2(n3538),
	.A3(n3537),
	.A4(n3536),
	.ZN(n3556));
   AOI22_X1 U4093 (.A1(REGISTERS[94]),
	.A2(FE_OFN131_n3570),
	.B1(REGISTERS[30]),
	.B2(FE_OFN108_n3569),
	.ZN(n3543));
   AOI22_X1 U4094 (.A1(REGISTERS[222]),
	.A2(FE_OFN46_n3572),
	.B1(REGISTERS[158]),
	.B2(FE_OFN7_n3571),
	.ZN(n3542));
   AOI22_X1 U4095 (.A1(REGISTERS[126]),
	.A2(FE_OFN3_n3574),
	.B1(REGISTERS[62]),
	.B2(FE_OFN133_n3573),
	.ZN(n3541));
   AOI22_X1 U4096 (.A1(REGISTERS[254]),
	.A2(FE_OFN105_n3576),
	.B1(REGISTERS[190]),
	.B2(FE_OFN49_n3575),
	.ZN(n3540));
   AND4_X1 U4097 (.A1(n3543),
	.A2(n3542),
	.A3(n3541),
	.A4(n3540),
	.ZN(n3555));
   AOI22_X1 U4098 (.A1(REGISTERS[862]),
	.A2(FE_OFN132_n3570),
	.B1(REGISTERS[798]),
	.B2(FE_OFN109_n3569),
	.ZN(n3547));
   AOI22_X1 U4099 (.A1(REGISTERS[990]),
	.A2(FE_OFN47_n3572),
	.B1(REGISTERS[926]),
	.B2(FE_OFN7_n3571),
	.ZN(n3546));
   AOI22_X1 U4100 (.A1(REGISTERS[894]),
	.A2(FE_OFN5_n3574),
	.B1(REGISTERS[830]),
	.B2(FE_OFN134_n3573),
	.ZN(n3545));
   AOI22_X1 U4101 (.A1(REGISTERS[1022]),
	.A2(FE_OFN105_n3576),
	.B1(REGISTERS[958]),
	.B2(FE_OFN49_n3575),
	.ZN(n3544));
   NAND4_X1 U4102 (.A1(n3547),
	.A2(n3546),
	.A3(n3545),
	.A4(n3544),
	.ZN(n3553));
   AOI22_X1 U4103 (.A1(REGISTERS[606]),
	.A2(FE_OFN132_n3570),
	.B1(REGISTERS[542]),
	.B2(FE_OFN109_n3569),
	.ZN(n3551));
   AOI22_X1 U4104 (.A1(REGISTERS[734]),
	.A2(FE_OFN47_n3572),
	.B1(REGISTERS[670]),
	.B2(FE_OFN7_n3571),
	.ZN(n3550));
   AOI22_X1 U4105 (.A1(REGISTERS[638]),
	.A2(FE_OFN5_n3574),
	.B1(REGISTERS[574]),
	.B2(FE_OFN134_n3573),
	.ZN(n3549));
   AOI22_X1 U4106 (.A1(REGISTERS[766]),
	.A2(FE_OFN105_n3576),
	.B1(REGISTERS[702]),
	.B2(FE_OFN49_n3575),
	.ZN(n3548));
   NAND4_X1 U4107 (.A1(n3551),
	.A2(n3550),
	.A3(n3549),
	.A4(n3548),
	.ZN(n3552));
   AOI22_X1 U4108 (.A1(n3553),
	.A2(FE_OFN33_n3584),
	.B1(n3552),
	.B2(FE_OFN31_n3582),
	.ZN(n3554));
   OAI221_X1 U4109 (.A(n3554),
	.B1(FE_OFN38_n3588),
	.B2(n3556),
	.C1(n3586),
	.C2(n3555),
	.ZN(N97));
   AOI22_X1 U4110 (.A1(REGISTERS[351]),
	.A2(FE_OFN131_n3570),
	.B1(REGISTERS[287]),
	.B2(FE_OFN108_n3569),
	.ZN(n3560));
   AOI22_X1 U4111 (.A1(REGISTERS[479]),
	.A2(n3572),
	.B1(REGISTERS[415]),
	.B2(n3571),
	.ZN(n3559));
   AOI22_X1 U4112 (.A1(REGISTERS[383]),
	.A2(n3574),
	.B1(REGISTERS[319]),
	.B2(n3573),
	.ZN(n3558));
   AOI22_X1 U4113 (.A1(REGISTERS[511]),
	.A2(FE_OFN106_n3576),
	.B1(REGISTERS[447]),
	.B2(FE_OFN48_n3575),
	.ZN(n3557));
   AND4_X1 U4114 (.A1(n3560),
	.A2(n3559),
	.A3(n3558),
	.A4(n3557),
	.ZN(n3589));
   AOI22_X1 U4115 (.A1(REGISTERS[95]),
	.A2(FE_OFN131_n3570),
	.B1(REGISTERS[31]),
	.B2(FE_OFN108_n3569),
	.ZN(n3564));
   AOI22_X1 U4116 (.A1(REGISTERS[223]),
	.A2(n3572),
	.B1(REGISTERS[159]),
	.B2(n3571),
	.ZN(n3563));
   AOI22_X1 U4117 (.A1(REGISTERS[127]),
	.A2(n3574),
	.B1(REGISTERS[63]),
	.B2(n3573),
	.ZN(n3562));
   AOI22_X1 U4118 (.A1(REGISTERS[255]),
	.A2(FE_OFN106_n3576),
	.B1(REGISTERS[191]),
	.B2(FE_OFN48_n3575),
	.ZN(n3561));
   AND4_X1 U4119 (.A1(n3564),
	.A2(n3563),
	.A3(n3562),
	.A4(n3561),
	.ZN(n3587));
   AOI22_X1 U4120 (.A1(REGISTERS[863]),
	.A2(FE_OFN131_n3570),
	.B1(REGISTERS[799]),
	.B2(FE_OFN108_n3569),
	.ZN(n3568));
   AOI22_X1 U4121 (.A1(REGISTERS[991]),
	.A2(FE_OFN46_n3572),
	.B1(REGISTERS[927]),
	.B2(n3571),
	.ZN(n3567));
   AOI22_X1 U4122 (.A1(REGISTERS[895]),
	.A2(n3574),
	.B1(REGISTERS[831]),
	.B2(n3573),
	.ZN(n3566));
   AOI22_X1 U4123 (.A1(REGISTERS[1023]),
	.A2(FE_OFN106_n3576),
	.B1(REGISTERS[959]),
	.B2(FE_OFN48_n3575),
	.ZN(n3565));
   NAND4_X1 U4124 (.A1(n3568),
	.A2(n3567),
	.A3(n3566),
	.A4(n3565),
	.ZN(n3583));
   AOI22_X1 U4125 (.A1(REGISTERS[607]),
	.A2(FE_OFN131_n3570),
	.B1(REGISTERS[543]),
	.B2(FE_OFN108_n3569),
	.ZN(n3580));
   AOI22_X1 U4126 (.A1(REGISTERS[735]),
	.A2(FE_OFN46_n3572),
	.B1(REGISTERS[671]),
	.B2(n3571),
	.ZN(n3579));
   AOI22_X1 U4127 (.A1(REGISTERS[639]),
	.A2(n3574),
	.B1(REGISTERS[575]),
	.B2(n3573),
	.ZN(n3578));
   AOI22_X1 U4128 (.A1(REGISTERS[767]),
	.A2(FE_OFN106_n3576),
	.B1(REGISTERS[703]),
	.B2(FE_OFN48_n3575),
	.ZN(n3577));
   NAND4_X1 U4129 (.A1(n3580),
	.A2(n3579),
	.A3(n3578),
	.A4(n3577),
	.ZN(n3581));
   AOI22_X1 U4130 (.A1(FE_OFN33_n3584),
	.A2(n3583),
	.B1(FE_OFN31_n3582),
	.B2(n3581),
	.ZN(n3585));
   OAI221_X1 U4131 (.A(n3585),
	.B1(n3589),
	.B2(FE_OFN38_n3588),
	.C1(n3587),
	.C2(n3586),
	.ZN(N96));
   INV_X1 U4140 (.A(ADD_WR[0]),
	.ZN(n4040));
endmodule

module decode_unit_DW01_add_0 (
	A, 
	B, 
	CI, 
	SUM, 
	CO);
   input [31:0] A;
   input [31:0] B;
   input CI;
   output [31:0] SUM;
   output CO;

   // Internal wires
   wire n2;
   wire n9;
   wire n16;
   wire n17;
   wire n18;
   wire n19;
   wire n20;
   wire n21;
   wire n22;
   wire n23;
   wire n28;
   wire n31;
   wire n35;
   wire n36;
   wire n37;
   wire n38;
   wire n39;
   wire n40;
   wire n41;
   wire n42;
   wire n43;
   wire n44;
   wire n45;
   wire n46;
   wire n47;
   wire n48;
   wire n49;
   wire n50;
   wire n51;
   wire n52;
   wire n53;
   wire n54;
   wire n55;
   wire n57;
   wire n58;
   wire n59;
   wire n60;
   wire n61;
   wire n62;
   wire n63;
   wire n64;
   wire n65;
   wire n66;
   wire n67;
   wire n68;
   wire n69;
   wire n70;
   wire n71;
   wire n72;
   wire n73;
   wire n74;
   wire n75;
   wire n76;
   wire n78;
   wire n80;
   wire n81;
   wire n82;
   wire n83;
   wire n84;
   wire n85;
   wire n86;
   wire n87;
   wire n88;
   wire n89;
   wire n90;
   wire n91;
   wire n92;
   wire n93;
   wire n94;
   wire n95;
   wire n102;
   wire n104;
   wire n105;
   wire n106;
   wire n107;
   wire n108;
   wire n109;
   wire n110;
   wire n111;
   wire n112;
   wire n113;
   wire n114;
   wire n115;
   wire n118;
   wire n119;
   wire n120;
   wire n121;
   wire n122;
   wire n123;
   wire n124;
   wire n125;
   wire n126;
   wire n127;
   wire n128;
   wire n129;
   wire n130;
   wire n131;
   wire n132;
   wire n133;
   wire n134;
   wire n135;
   wire n136;
   wire n137;
   wire n138;
   wire n139;
   wire n140;
   wire n141;
   wire n142;
   wire n143;
   wire n144;
   wire n145;
   wire n147;
   wire [31:2] carry;

   FA_X1 U1_22 (.A(A[22]),
	.B(B[22]),
	.CI(carry[22]),
	.CO(carry[23]),
	.S(SUM[22]));
   FA_X1 U1_16 (.A(A[16]),
	.B(B[16]),
	.CI(carry[16]),
	.CO(carry[17]),
	.S(SUM[16]));
   FA_X1 U1_6 (.A(A[6]),
	.B(B[6]),
	.CI(carry[6]),
	.CO(carry[7]),
	.S(SUM[6]));
   FA_X1 U1_1 (.A(n147),
	.B(A[1]),
	.CI(B[1]),
	.CO(carry[2]),
	.S(SUM[1]));
   XNOR2_X1 U2 (.A(B[31]),
	.B(A[31]),
	.ZN(n2));
   NAND3_X1 U9 (.A1(n111),
	.A2(n110),
	.A3(n109),
	.ZN(n9));
   XOR2_X1 U16 (.A(B[11]),
	.B(A[11]),
	.Z(n16));
   XOR2_X1 U17 (.A(n9),
	.B(n16),
	.Z(SUM[11]));
   NAND2_X1 U18 (.A1(n9),
	.A2(B[11]),
	.ZN(n17));
   NAND2_X1 U19 (.A1(n9),
	.A2(A[11]),
	.ZN(n18));
   NAND2_X1 U20 (.A1(B[11]),
	.A2(A[11]),
	.ZN(n19));
   NAND3_X1 U21 (.A1(n17),
	.A2(n18),
	.A3(n19),
	.ZN(carry[12]));
   XOR2_X1 U22 (.A(B[17]),
	.B(A[17]),
	.Z(n20));
   XOR2_X1 U23 (.A(carry[17]),
	.B(n20),
	.Z(SUM[17]));
   NAND2_X1 U24 (.A1(carry[17]),
	.A2(B[17]),
	.ZN(n21));
   NAND2_X1 U25 (.A1(carry[17]),
	.A2(A[17]),
	.ZN(n22));
   NAND2_X1 U26 (.A1(B[17]),
	.A2(A[17]),
	.ZN(n23));
   NAND3_X1 U27 (.A1(n21),
	.A2(n22),
	.A3(n23),
	.ZN(carry[18]));
   NAND3_X1 U32 (.A1(n119),
	.A2(n120),
	.A3(n121),
	.ZN(n28));
   NAND3_X1 U35 (.A1(n141),
	.A2(n140),
	.A3(n139),
	.ZN(n31));
   XOR2_X1 U39 (.A(B[30]),
	.B(A[30]),
	.Z(n35));
   XOR2_X1 U40 (.A(n28),
	.B(n35),
	.Z(SUM[30]));
   NAND2_X1 U41 (.A1(n28),
	.A2(B[30]),
	.ZN(n36));
   NAND2_X1 U42 (.A1(n28),
	.A2(A[30]),
	.ZN(n37));
   NAND2_X1 U43 (.A1(B[30]),
	.A2(A[30]),
	.ZN(n38));
   NAND3_X1 U44 (.A1(n36),
	.A2(n37),
	.A3(n38),
	.ZN(carry[31]));
   XOR2_X1 U45 (.A(B[15]),
	.B(A[15]),
	.Z(n39));
   XOR2_X1 U46 (.A(n31),
	.B(n39),
	.Z(SUM[15]));
   NAND2_X1 U47 (.A1(n31),
	.A2(B[15]),
	.ZN(n40));
   NAND2_X1 U48 (.A1(n31),
	.A2(A[15]),
	.ZN(n41));
   NAND2_X1 U49 (.A1(B[15]),
	.A2(A[15]),
	.ZN(n42));
   NAND3_X1 U50 (.A1(n40),
	.A2(n41),
	.A3(n42),
	.ZN(carry[16]));
   XNOR2_X1 U51 (.A(carry[31]),
	.B(n2),
	.ZN(SUM[31]));
   XOR2_X1 U52 (.A(A[18]),
	.B(B[18]),
	.Z(n43));
   XOR2_X1 U53 (.A(n43),
	.B(carry[18]),
	.Z(SUM[18]));
   NAND2_X1 U54 (.A1(A[18]),
	.A2(B[18]),
	.ZN(n44));
   NAND2_X1 U55 (.A1(A[18]),
	.A2(carry[18]),
	.ZN(n45));
   NAND2_X1 U56 (.A1(B[18]),
	.A2(carry[18]),
	.ZN(n46));
   NAND3_X1 U57 (.A1(n44),
	.A2(n45),
	.A3(n46),
	.ZN(carry[19]));
   XOR2_X1 U58 (.A(A[19]),
	.B(B[19]),
	.Z(n47));
   XOR2_X1 U59 (.A(n47),
	.B(carry[19]),
	.Z(SUM[19]));
   NAND2_X1 U60 (.A1(A[19]),
	.A2(B[19]),
	.ZN(n48));
   NAND2_X1 U61 (.A1(A[19]),
	.A2(carry[19]),
	.ZN(n49));
   NAND2_X1 U62 (.A1(B[19]),
	.A2(carry[19]),
	.ZN(n50));
   NAND3_X1 U63 (.A1(n48),
	.A2(n49),
	.A3(n50),
	.ZN(carry[20]));
   XOR2_X1 U64 (.A(B[26]),
	.B(A[26]),
	.Z(n51));
   XOR2_X1 U65 (.A(carry[26]),
	.B(n51),
	.Z(SUM[26]));
   NAND2_X1 U66 (.A1(carry[26]),
	.A2(B[26]),
	.ZN(n52));
   NAND2_X1 U67 (.A1(carry[26]),
	.A2(A[26]),
	.ZN(n53));
   NAND2_X1 U68 (.A1(B[26]),
	.A2(A[26]),
	.ZN(n54));
   NAND3_X1 U69 (.A1(n52),
	.A2(n53),
	.A3(n54),
	.ZN(carry[27]));
   NAND3_X1 U70 (.A1(n144),
	.A2(n143),
	.A3(n145),
	.ZN(n55));
   XOR2_X1 U72 (.A(B[25]),
	.B(A[25]),
	.Z(n57));
   XOR2_X1 U73 (.A(carry[25]),
	.B(n57),
	.Z(SUM[25]));
   NAND2_X1 U74 (.A1(carry[25]),
	.A2(B[25]),
	.ZN(n58));
   NAND2_X1 U75 (.A1(carry[25]),
	.A2(A[25]),
	.ZN(n59));
   NAND2_X1 U76 (.A1(B[25]),
	.A2(A[25]),
	.ZN(n60));
   NAND3_X1 U77 (.A1(n58),
	.A2(n59),
	.A3(n60),
	.ZN(carry[26]));
   XOR2_X1 U78 (.A(B[20]),
	.B(A[20]),
	.Z(n61));
   XOR2_X1 U79 (.A(carry[20]),
	.B(n61),
	.Z(SUM[20]));
   NAND2_X1 U80 (.A1(carry[20]),
	.A2(B[20]),
	.ZN(n62));
   NAND2_X1 U81 (.A1(carry[20]),
	.A2(A[20]),
	.ZN(n63));
   NAND2_X1 U82 (.A1(B[20]),
	.A2(A[20]),
	.ZN(n64));
   NAND3_X1 U83 (.A1(n62),
	.A2(n63),
	.A3(n64),
	.ZN(carry[21]));
   XOR2_X1 U84 (.A(B[4]),
	.B(A[4]),
	.Z(n65));
   XOR2_X1 U85 (.A(n55),
	.B(n65),
	.Z(SUM[4]));
   NAND2_X1 U86 (.A1(n55),
	.A2(B[4]),
	.ZN(n66));
   NAND2_X1 U87 (.A1(n55),
	.A2(A[4]),
	.ZN(n67));
   NAND2_X1 U88 (.A1(B[4]),
	.A2(A[4]),
	.ZN(n68));
   NAND3_X1 U89 (.A1(n67),
	.A2(n66),
	.A3(n68),
	.ZN(carry[5]));
   XOR2_X1 U90 (.A(B[21]),
	.B(A[21]),
	.Z(n69));
   XOR2_X1 U91 (.A(carry[21]),
	.B(n69),
	.Z(SUM[21]));
   NAND2_X1 U92 (.A1(carry[21]),
	.A2(B[21]),
	.ZN(n70));
   NAND2_X1 U93 (.A1(carry[21]),
	.A2(A[21]),
	.ZN(n71));
   NAND2_X1 U94 (.A1(B[21]),
	.A2(A[21]),
	.ZN(n72));
   NAND3_X1 U95 (.A1(n70),
	.A2(n71),
	.A3(n72),
	.ZN(carry[22]));
   XOR2_X1 U96 (.A(B[5]),
	.B(A[5]),
	.Z(n73));
   XOR2_X1 U97 (.A(carry[5]),
	.B(n73),
	.Z(SUM[5]));
   NAND2_X1 U98 (.A1(carry[5]),
	.A2(B[5]),
	.ZN(n74));
   NAND2_X1 U99 (.A1(carry[5]),
	.A2(A[5]),
	.ZN(n75));
   NAND2_X1 U100 (.A1(B[5]),
	.A2(A[5]),
	.ZN(n76));
   NAND3_X1 U101 (.A1(n74),
	.A2(n75),
	.A3(n76),
	.ZN(carry[6]));
   NAND3_X1 U103 (.A1(n90),
	.A2(n89),
	.A3(n91),
	.ZN(n78));
   XOR2_X1 U105 (.A(B[23]),
	.B(A[23]),
	.Z(n80));
   XOR2_X1 U106 (.A(carry[23]),
	.B(n80),
	.Z(SUM[23]));
   NAND2_X1 U107 (.A1(carry[23]),
	.A2(B[23]),
	.ZN(n81));
   NAND2_X1 U108 (.A1(carry[23]),
	.A2(A[23]),
	.ZN(n82));
   NAND2_X1 U109 (.A1(B[23]),
	.A2(A[23]),
	.ZN(n83));
   NAND3_X1 U110 (.A1(n81),
	.A2(n82),
	.A3(n83),
	.ZN(carry[24]));
   XOR2_X1 U111 (.A(B[27]),
	.B(A[27]),
	.Z(n84));
   XOR2_X1 U112 (.A(carry[27]),
	.B(n84),
	.Z(SUM[27]));
   NAND2_X1 U113 (.A1(carry[27]),
	.A2(B[27]),
	.ZN(n85));
   NAND2_X1 U114 (.A1(carry[27]),
	.A2(A[27]),
	.ZN(n86));
   NAND2_X1 U115 (.A1(B[27]),
	.A2(A[27]),
	.ZN(n87));
   NAND3_X1 U116 (.A1(n85),
	.A2(n86),
	.A3(n87),
	.ZN(carry[28]));
   XOR2_X1 U117 (.A(B[2]),
	.B(A[2]),
	.Z(n88));
   XOR2_X1 U118 (.A(carry[2]),
	.B(n88),
	.Z(SUM[2]));
   NAND2_X1 U119 (.A1(carry[2]),
	.A2(B[2]),
	.ZN(n89));
   NAND2_X1 U120 (.A1(carry[2]),
	.A2(A[2]),
	.ZN(n90));
   NAND2_X1 U121 (.A1(B[2]),
	.A2(A[2]),
	.ZN(n91));
   NAND3_X1 U122 (.A1(n89),
	.A2(n90),
	.A3(n91),
	.ZN(carry[3]));
   XOR2_X1 U123 (.A(B[12]),
	.B(A[12]),
	.Z(n92));
   XOR2_X1 U124 (.A(carry[12]),
	.B(n92),
	.Z(SUM[12]));
   NAND2_X1 U125 (.A1(carry[12]),
	.A2(B[12]),
	.ZN(n93));
   NAND2_X1 U126 (.A1(carry[12]),
	.A2(A[12]),
	.ZN(n94));
   NAND2_X1 U127 (.A1(B[12]),
	.A2(A[12]),
	.ZN(n95));
   NAND3_X1 U128 (.A1(n93),
	.A2(n94),
	.A3(n95),
	.ZN(carry[13]));
   NAND3_X1 U135 (.A1(n107),
	.A2(n106),
	.A3(n105),
	.ZN(n102));
   XOR2_X1 U137 (.A(A[9]),
	.B(B[9]),
	.Z(n104));
   XOR2_X1 U138 (.A(n104),
	.B(carry[9]),
	.Z(SUM[9]));
   NAND2_X1 U139 (.A1(A[9]),
	.A2(B[9]),
	.ZN(n105));
   NAND2_X1 U140 (.A1(A[9]),
	.A2(carry[9]),
	.ZN(n106));
   NAND2_X1 U141 (.A1(B[9]),
	.A2(carry[9]),
	.ZN(n107));
   NAND3_X1 U142 (.A1(n105),
	.A2(n106),
	.A3(n107),
	.ZN(carry[10]));
   XOR2_X1 U143 (.A(A[10]),
	.B(B[10]),
	.Z(n108));
   XOR2_X1 U144 (.A(n108),
	.B(carry[10]),
	.Z(SUM[10]));
   NAND2_X1 U145 (.A1(A[10]),
	.A2(B[10]),
	.ZN(n109));
   NAND2_X1 U146 (.A1(A[10]),
	.A2(n102),
	.ZN(n110));
   NAND2_X1 U147 (.A1(B[10]),
	.A2(carry[10]),
	.ZN(n111));
   XOR2_X1 U149 (.A(B[28]),
	.B(A[28]),
	.Z(n112));
   XOR2_X1 U150 (.A(carry[28]),
	.B(n112),
	.Z(SUM[28]));
   NAND2_X1 U151 (.A1(carry[28]),
	.A2(B[28]),
	.ZN(n113));
   NAND2_X1 U152 (.A1(carry[28]),
	.A2(A[28]),
	.ZN(n114));
   NAND2_X1 U153 (.A1(B[28]),
	.A2(A[28]),
	.ZN(n115));
   NAND3_X1 U154 (.A1(n113),
	.A2(n114),
	.A3(n115),
	.ZN(carry[29]));
   XOR2_X1 U157 (.A(B[29]),
	.B(A[29]),
	.Z(n118));
   XOR2_X1 U158 (.A(carry[29]),
	.B(n118),
	.Z(SUM[29]));
   NAND2_X1 U159 (.A1(carry[29]),
	.A2(B[29]),
	.ZN(n119));
   NAND2_X1 U160 (.A1(carry[29]),
	.A2(A[29]),
	.ZN(n120));
   NAND2_X1 U161 (.A1(B[29]),
	.A2(A[29]),
	.ZN(n121));
   XOR2_X1 U163 (.A(A[7]),
	.B(B[7]),
	.Z(n122));
   XOR2_X1 U164 (.A(n122),
	.B(carry[7]),
	.Z(SUM[7]));
   NAND2_X1 U165 (.A1(A[7]),
	.A2(B[7]),
	.ZN(n123));
   NAND2_X1 U166 (.A1(A[7]),
	.A2(carry[7]),
	.ZN(n124));
   NAND2_X1 U167 (.A1(B[7]),
	.A2(carry[7]),
	.ZN(n125));
   NAND3_X1 U168 (.A1(n123),
	.A2(n124),
	.A3(n125),
	.ZN(carry[8]));
   XOR2_X1 U169 (.A(A[8]),
	.B(B[8]),
	.Z(n126));
   XOR2_X1 U170 (.A(n126),
	.B(carry[8]),
	.Z(SUM[8]));
   NAND2_X1 U171 (.A1(A[8]),
	.A2(B[8]),
	.ZN(n127));
   NAND2_X1 U172 (.A1(A[8]),
	.A2(carry[8]),
	.ZN(n128));
   NAND2_X1 U173 (.A1(carry[8]),
	.A2(B[8]),
	.ZN(n129));
   NAND3_X1 U174 (.A1(n127),
	.A2(n128),
	.A3(n129),
	.ZN(carry[9]));
   XOR2_X1 U175 (.A(B[24]),
	.B(A[24]),
	.Z(n130));
   XOR2_X1 U176 (.A(carry[24]),
	.B(n130),
	.Z(SUM[24]));
   NAND2_X1 U177 (.A1(carry[24]),
	.A2(B[24]),
	.ZN(n131));
   NAND2_X1 U178 (.A1(carry[24]),
	.A2(A[24]),
	.ZN(n132));
   NAND2_X1 U179 (.A1(B[24]),
	.A2(A[24]),
	.ZN(n133));
   NAND3_X1 U180 (.A1(n131),
	.A2(n132),
	.A3(n133),
	.ZN(carry[25]));
   XOR2_X1 U181 (.A(A[13]),
	.B(B[13]),
	.Z(n134));
   XOR2_X1 U182 (.A(n134),
	.B(carry[13]),
	.Z(SUM[13]));
   NAND2_X1 U183 (.A1(A[13]),
	.A2(B[13]),
	.ZN(n135));
   NAND2_X1 U184 (.A1(carry[13]),
	.A2(A[13]),
	.ZN(n136));
   NAND2_X1 U185 (.A1(carry[13]),
	.A2(B[13]),
	.ZN(n137));
   NAND3_X1 U186 (.A1(n135),
	.A2(n136),
	.A3(n137),
	.ZN(carry[14]));
   XOR2_X1 U187 (.A(A[14]),
	.B(B[14]),
	.Z(n138));
   XOR2_X1 U188 (.A(n138),
	.B(carry[14]),
	.Z(SUM[14]));
   NAND2_X1 U189 (.A1(A[14]),
	.A2(B[14]),
	.ZN(n139));
   NAND2_X1 U190 (.A1(carry[14]),
	.A2(A[14]),
	.ZN(n140));
   NAND2_X1 U191 (.A1(B[14]),
	.A2(carry[14]),
	.ZN(n141));
   XOR2_X1 U193 (.A(B[3]),
	.B(A[3]),
	.Z(n142));
   XOR2_X1 U194 (.A(carry[3]),
	.B(n142),
	.Z(SUM[3]));
   NAND2_X1 U195 (.A1(n78),
	.A2(B[3]),
	.ZN(n143));
   NAND2_X1 U196 (.A1(carry[3]),
	.A2(A[3]),
	.ZN(n144));
   NAND2_X1 U197 (.A1(B[3]),
	.A2(A[3]),
	.ZN(n145));
   XOR2_X1 U199 (.A(B[0]),
	.B(A[0]),
	.Z(SUM[0]));
   AND2_X1 U200 (.A1(B[0]),
	.A2(A[0]),
	.ZN(n147));
endmodule

module decode_unit (
	clk, 
	rst, 
	en, 
	RF_RD1, 
	RF_RD2, 
	RF_WR, 
	IF_FLUSH, 
	PC_IN, 
	IR_IN, 
	EXE_MEM_IN, 
	ADD_WR, 
	DATAIN, 
	MUX_IMM_SEL, 
	RF_OUT1_SEL, 
	RF_OUT2_SEL, 
	OPCODE, 
	FUNC3, 
	EQU_FLAG, 
	RF_OUT1, 
	RF_OUT2, 
	PC_OUT, 
	IMM, 
	JMP_ADDR, 
	RD, 
	RS1, 
	RS2);
   input clk;
   input rst;
   input en;
   input RF_RD1;
   input RF_RD2;
   input RF_WR;
   input IF_FLUSH;
   input [31:0] PC_IN;
   input [31:0] IR_IN;
   input [31:0] EXE_MEM_IN;
   input [4:0] ADD_WR;
   input [31:0] DATAIN;
   input [2:0] MUX_IMM_SEL;
   input [1:0] RF_OUT1_SEL;
   input [1:0] RF_OUT2_SEL;
   output [6:0] OPCODE;
   output [2:0] FUNC3;
   output EQU_FLAG;
   output [31:0] RF_OUT1;
   output [31:0] RF_OUT2;
   output [31:0] PC_OUT;
   output [31:0] IMM;
   output [31:0] JMP_ADDR;
   output [4:0] RD;
   output [4:0] RS1;
   output [4:0] RS2;

   // Internal wires
   wire FE_OFN93_n204;
   wire FE_OFN92_n170;
   wire FE_OFN35_n205;
   wire FE_OFN29_n171;
   wire FE_DBTN2_n10;
   wire FE_DBTN1_n11;
   wire n41;
   wire n43;
   wire n45;
   wire n47;
   wire n49;
   wire n51;
   wire n53;
   wire n55;
   wire n57;
   wire n59;
   wire n61;
   wire n63;
   wire n65;
   wire n67;
   wire n69;
   wire n71;
   wire n73;
   wire n75;
   wire n77;
   wire n79;
   wire n81;
   wire n83;
   wire n85;
   wire n87;
   wire n169;
   wire n170;
   wire n171;
   wire n172;
   wire n173;
   wire n174;
   wire n175;
   wire n176;
   wire n177;
   wire n178;
   wire n179;
   wire n180;
   wire n181;
   wire n182;
   wire n183;
   wire n184;
   wire n185;
   wire n186;
   wire n187;
   wire n188;
   wire n189;
   wire n190;
   wire n191;
   wire n192;
   wire n193;
   wire n194;
   wire n195;
   wire n196;
   wire n197;
   wire n198;
   wire n199;
   wire n200;
   wire n201;
   wire n202;
   wire n203;
   wire n204;
   wire n205;
   wire n206;
   wire n207;
   wire n208;
   wire n209;
   wire n210;
   wire n211;
   wire n212;
   wire n213;
   wire n214;
   wire n215;
   wire n216;
   wire n217;
   wire n218;
   wire n219;
   wire n220;
   wire n221;
   wire n222;
   wire n223;
   wire n224;
   wire n225;
   wire n226;
   wire n227;
   wire n228;
   wire n229;
   wire n230;
   wire n231;
   wire n232;
   wire n233;
   wire n234;
   wire n235;
   wire n236;
   wire n237;
   wire n238;
   wire n239;
   wire n240;
   wire n241;
   wire n242;
   wire n243;
   wire n244;
   wire n245;
   wire n246;
   wire n247;
   wire n248;
   wire n249;
   wire n251;
   wire n252;
   wire n253;
   wire n255;
   wire n256;
   wire n257;
   wire n258;
   wire n259;
   wire n260;
   wire n261;
   wire n262;
   wire n263;
   wire n264;
   wire n265;
   wire n266;
   wire n267;
   wire n268;
   wire n269;
   wire n270;
   wire n271;
   wire n272;
   wire n273;
   wire n274;
   wire n275;
   wire n276;
   wire n277;
   wire n278;
   wire n279;
   wire n280;
   wire n281;
   wire n282;
   wire n283;
   wire n284;
   wire n285;
   wire n286;
   wire n287;
   wire n288;
   wire n289;
   wire n290;
   wire n291;
   wire n292;
   wire n293;
   wire n294;
   wire n295;
   wire n296;
   wire n297;
   wire n298;
   wire n299;
   wire n300;
   wire n301;
   wire n302;
   wire n303;
   wire n304;
   wire n305;
   wire n306;
   wire n307;
   wire n308;
   wire n309;
   wire n310;
   wire n311;
   wire n312;
   wire n313;
   wire n314;
   wire n315;
   wire n316;
   wire n317;
   wire n318;
   wire n319;
   wire n320;
   wire n321;
   wire n322;
   wire n323;
   wire n324;
   wire n325;
   wire n326;
   wire n327;
   wire n328;
   wire n329;
   wire n330;
   wire n331;
   wire n332;
   wire n333;
   wire n334;
   wire n335;
   wire n336;
   wire n337;
   wire n338;
   wire n339;
   wire n340;
   wire n341;
   wire n342;
   wire n343;
   wire n344;
   wire n345;
   wire n346;
   wire n347;
   wire n348;
   wire n349;
   wire n350;
   wire n351;
   wire n352;
   wire n353;
   wire n354;
   wire n355;
   wire n356;
   wire n357;
   wire n358;
   wire n359;
   wire n4;
   wire n6;
   wire n7;
   wire n8;
   wire n9;
   wire n10;
   wire n11;
   wire n40;
   wire n42;
   wire n44;
   wire n46;
   wire n48;
   wire n50;
   wire n52;
   wire n54;
   wire n56;
   wire n58;
   wire n60;
   wire n62;
   wire n64;
   wire n66;
   wire n68;
   wire n70;
   wire n72;
   wire n74;
   wire n76;
   wire n78;
   wire n80;
   wire n82;
   wire n84;
   wire n86;
   wire n88;
   wire n89;
   wire n90;
   wire n91;
   wire n92;
   wire n93;
   wire n94;
   wire n95;
   wire n96;
   wire n97;
   wire n98;
   wire n99;
   wire n100;
   wire n101;
   wire n102;
   wire n103;
   wire n104;
   wire n105;
   wire n106;
   wire n107;
   wire n108;
   wire n109;
   wire n110;
   wire n111;
   wire n112;
   wire n113;
   wire n114;
   wire n115;
   wire n116;
   wire n117;
   wire n118;
   wire n119;
   wire n120;
   wire n121;
   wire n122;
   wire n123;
   wire n124;
   wire n125;
   wire n126;
   wire n127;
   wire n128;
   wire n129;
   wire n130;
   wire n131;
   wire n132;
   wire n133;
   wire n134;
   wire n135;
   wire n136;
   wire n137;
   wire n138;
   wire n139;
   wire n140;
   wire n141;
   wire n142;
   wire n143;
   wire n144;
   wire n145;
   wire n146;
   wire n147;
   wire n148;
   wire n149;
   wire n150;
   wire n151;
   wire n152;
   wire n153;
   wire n154;
   wire n155;
   wire n156;
   wire n157;
   wire n158;
   wire n159;
   wire n160;
   wire n161;
   wire n162;
   wire n163;
   wire n164;
   wire n165;
   wire n166;
   wire n167;
   wire n168;
   wire n250;
   wire n254;
   wire n360;
   wire n361;
   wire n362;
   wire n363;
   wire n364;
   wire n365;
   wire n366;
   wire n367;
   wire n368;
   wire n369;
   wire n370;
   wire n371;
   wire n372;
   wire n373;
   wire n374;
   wire n375;
   wire n376;
   wire n377;
   wire n378;
   wire n379;
   wire n380;
   wire n381;
   wire n382;
   wire n383;
   wire n384;
   wire n385;
   wire [30:25] currIR;
   wire [31:0] RF_OUT1_m;
   wire [31:0] RF_OUT2_m;

   BUF_X2 FE_OFC93_n204 (.A(n204),
	.Z(FE_OFN93_n204));
   BUF_X2 FE_OFC92_n170 (.A(n170),
	.Z(FE_OFN92_n170));
   BUF_X2 FE_OFC35_n205 (.A(n205),
	.Z(FE_OFN35_n205));
   BUF_X2 FE_OFC29_n171 (.A(n171),
	.Z(FE_OFN29_n171));
   INV_X2 FE_DBTC2_n10 (.A(n10),
	.ZN(FE_DBTN2_n10));
   INV_X2 FE_DBTC1_n11 (.A(n11),
	.ZN(FE_DBTN1_n11));
   DFF_X1 currPC_reg_31_ (.D(n130),
	.CK(clk),
	.Q(PC_OUT[31]));
   DFF_X1 currPC_reg_30_ (.D(n131),
	.CK(clk),
	.Q(PC_OUT[30]));
   DFF_X1 currPC_reg_29_ (.D(n132),
	.CK(clk),
	.Q(PC_OUT[29]));
   DFF_X1 currPC_reg_28_ (.D(n133),
	.CK(clk),
	.Q(PC_OUT[28]));
   DFF_X1 currPC_reg_27_ (.D(n134),
	.CK(clk),
	.Q(PC_OUT[27]));
   DFF_X1 currPC_reg_26_ (.D(n135),
	.CK(clk),
	.Q(PC_OUT[26]));
   DFF_X1 currPC_reg_25_ (.D(n136),
	.CK(clk),
	.Q(PC_OUT[25]));
   DFF_X1 currPC_reg_24_ (.D(n137),
	.CK(clk),
	.Q(PC_OUT[24]));
   DFF_X1 currPC_reg_23_ (.D(n138),
	.CK(clk),
	.Q(PC_OUT[23]));
   DFF_X1 currPC_reg_22_ (.D(n139),
	.CK(clk),
	.Q(PC_OUT[22]));
   DFF_X1 currPC_reg_21_ (.D(n140),
	.CK(clk),
	.Q(PC_OUT[21]));
   DFF_X1 currPC_reg_20_ (.D(n141),
	.CK(clk),
	.Q(PC_OUT[20]));
   DFF_X1 currPC_reg_19_ (.D(n142),
	.CK(clk),
	.Q(PC_OUT[19]));
   DFF_X1 currPC_reg_18_ (.D(n143),
	.CK(clk),
	.Q(PC_OUT[18]));
   DFF_X1 currPC_reg_17_ (.D(n144),
	.CK(clk),
	.Q(PC_OUT[17]));
   DFF_X1 currPC_reg_16_ (.D(n145),
	.CK(clk),
	.Q(PC_OUT[16]));
   DFF_X1 currPC_reg_15_ (.D(n146),
	.CK(clk),
	.Q(PC_OUT[15]));
   DFF_X1 currPC_reg_14_ (.D(n147),
	.CK(clk),
	.Q(PC_OUT[14]));
   DFF_X1 currPC_reg_13_ (.D(n148),
	.CK(clk),
	.Q(PC_OUT[13]));
   DFF_X1 currPC_reg_12_ (.D(n149),
	.CK(clk),
	.Q(PC_OUT[12]));
   DFF_X1 currPC_reg_11_ (.D(n150),
	.CK(clk),
	.Q(PC_OUT[11]));
   DFF_X1 currPC_reg_10_ (.D(n151),
	.CK(clk),
	.Q(PC_OUT[10]));
   DFF_X1 currPC_reg_9_ (.D(n152),
	.CK(clk),
	.Q(PC_OUT[9]));
   DFF_X1 currPC_reg_8_ (.D(n153),
	.CK(clk),
	.Q(PC_OUT[8]));
   DFF_X1 currPC_reg_7_ (.D(n154),
	.CK(clk),
	.Q(PC_OUT[7]));
   DFF_X1 currPC_reg_6_ (.D(n155),
	.CK(clk),
	.Q(PC_OUT[6]));
   DFF_X1 currPC_reg_5_ (.D(n156),
	.CK(clk),
	.Q(PC_OUT[5]));
   DFF_X1 currPC_reg_4_ (.D(n157),
	.CK(clk),
	.Q(PC_OUT[4]));
   DFF_X1 currPC_reg_3_ (.D(n158),
	.CK(clk),
	.Q(PC_OUT[3]));
   DFF_X1 currPC_reg_2_ (.D(n159),
	.CK(clk),
	.Q(PC_OUT[2]));
   DFF_X1 currPC_reg_1_ (.D(n160),
	.CK(clk),
	.Q(PC_OUT[1]));
   DFF_X1 currPC_reg_0_ (.D(n161),
	.CK(clk),
	.Q(PC_OUT[0]));
   DFF_X1 currIR_reg_31_ (.D(n40),
	.CK(clk),
	.Q(IMM[31]));
   DFF_X1 currIR_reg_30_ (.D(n42),
	.CK(clk),
	.Q(currIR[30]),
	.QN(n41));
   DFF_X1 currIR_reg_29_ (.D(n44),
	.CK(clk),
	.Q(currIR[29]),
	.QN(n43));
   DFF_X1 currIR_reg_28_ (.D(n46),
	.CK(clk),
	.Q(currIR[28]),
	.QN(n45));
   DFF_X1 currIR_reg_27_ (.D(n48),
	.CK(clk),
	.Q(currIR[27]),
	.QN(n47));
   DFF_X1 currIR_reg_26_ (.D(n50),
	.CK(clk),
	.Q(currIR[26]),
	.QN(n49));
   DFF_X1 currIR_reg_25_ (.D(n52),
	.CK(clk),
	.Q(currIR[25]),
	.QN(n51));
   DFF_X1 currIR_reg_24_ (.D(n54),
	.CK(clk),
	.Q(RS2[4]),
	.QN(n53));
   DFF_X1 currIR_reg_23_ (.D(n56),
	.CK(clk),
	.Q(RS2[3]),
	.QN(n55));
   DFF_X1 currIR_reg_22_ (.D(n58),
	.CK(clk),
	.Q(RS2[2]),
	.QN(n57));
   DFF_X1 currIR_reg_21_ (.D(n60),
	.CK(clk),
	.Q(RS2[1]),
	.QN(n59));
   DFF_X1 currIR_reg_20_ (.D(n62),
	.CK(clk),
	.Q(RS2[0]),
	.QN(n61));
   DFF_X1 currIR_reg_19_ (.D(n64),
	.CK(clk),
	.Q(RS1[4]),
	.QN(n63));
   DFF_X1 currIR_reg_18_ (.D(n66),
	.CK(clk),
	.Q(RS1[3]),
	.QN(n65));
   DFF_X1 currIR_reg_17_ (.D(n68),
	.CK(clk),
	.Q(RS1[2]),
	.QN(n67));
   DFF_X1 currIR_reg_16_ (.D(n70),
	.CK(clk),
	.Q(RS1[1]),
	.QN(n69));
   DFF_X1 currIR_reg_15_ (.D(n72),
	.CK(clk),
	.Q(RS1[0]),
	.QN(n71));
   DFF_X1 currIR_reg_14_ (.D(n74),
	.CK(clk),
	.Q(FUNC3[2]),
	.QN(n73));
   DFF_X1 currIR_reg_13_ (.D(n76),
	.CK(clk),
	.Q(FUNC3[1]),
	.QN(n75));
   DFF_X1 currIR_reg_12_ (.D(n78),
	.CK(clk),
	.Q(FUNC3[0]),
	.QN(n77));
   DFF_X1 currIR_reg_11_ (.D(n80),
	.CK(clk),
	.Q(RD[4]),
	.QN(n79));
   DFF_X1 currIR_reg_10_ (.D(n82),
	.CK(clk),
	.Q(RD[3]),
	.QN(n81));
   DFF_X1 currIR_reg_9_ (.D(n84),
	.CK(clk),
	.Q(RD[2]),
	.QN(n83));
   DFF_X1 currIR_reg_8_ (.D(n86),
	.CK(clk),
	.Q(RD[1]),
	.QN(n85));
   DFF_X1 currIR_reg_7_ (.D(n88),
	.CK(clk),
	.Q(RD[0]),
	.QN(n87));
   DFF_X1 currIR_reg_6_ (.D(n89),
	.CK(clk),
	.Q(OPCODE[6]));
   DFF_X1 currIR_reg_5_ (.D(n90),
	.CK(clk),
	.Q(OPCODE[5]));
   DFF_X1 currIR_reg_4_ (.D(n91),
	.CK(clk),
	.Q(OPCODE[4]));
   DFF_X1 currIR_reg_2_ (.D(n93),
	.CK(clk),
	.Q(OPCODE[2]));
   NAND2_X1 U252 (.A1(n351),
	.A2(n4),
	.ZN(n354));
   AND2_X1 U253 (.A1(n356),
	.A2(n9),
	.ZN(n351));
   XOR2_X1 U395 (.A(RF_OUT2[31]),
	.B(RF_OUT1[31]),
	.Z(n246));
   XOR2_X1 U396 (.A(RF_OUT2[30]),
	.B(RF_OUT1[30]),
	.Z(n245));
   XOR2_X1 U397 (.A(RF_OUT2[29]),
	.B(RF_OUT1[29]),
	.Z(n244));
   XOR2_X1 U398 (.A(RF_OUT2[28]),
	.B(RF_OUT1[28]),
	.Z(n243));
   XOR2_X1 U399 (.A(RF_OUT2[27]),
	.B(RF_OUT1[27]),
	.Z(n264));
   XOR2_X1 U400 (.A(RF_OUT2[26]),
	.B(RF_OUT1[26]),
	.Z(n263));
   XOR2_X1 U401 (.A(RF_OUT2[25]),
	.B(RF_OUT1[25]),
	.Z(n262));
   XOR2_X1 U402 (.A(RF_OUT2[24]),
	.B(RF_OUT1[24]),
	.Z(n261));
   XOR2_X1 U403 (.A(RF_OUT2[23]),
	.B(RF_OUT1[23]),
	.Z(n276));
   XOR2_X1 U404 (.A(RF_OUT2[22]),
	.B(RF_OUT1[22]),
	.Z(n275));
   XOR2_X1 U405 (.A(RF_OUT2[21]),
	.B(RF_OUT1[21]),
	.Z(n274));
   XOR2_X1 U406 (.A(RF_OUT2[20]),
	.B(RF_OUT1[20]),
	.Z(n273));
   XOR2_X1 U407 (.A(RF_OUT2[19]),
	.B(RF_OUT1[19]),
	.Z(n288));
   XOR2_X1 U408 (.A(RF_OUT2[18]),
	.B(RF_OUT1[18]),
	.Z(n287));
   XOR2_X1 U409 (.A(RF_OUT2[17]),
	.B(RF_OUT1[17]),
	.Z(n286));
   XOR2_X1 U410 (.A(RF_OUT2[16]),
	.B(RF_OUT1[16]),
	.Z(n285));
   XOR2_X1 U411 (.A(RF_OUT2[15]),
	.B(RF_OUT1[15]),
	.Z(n304));
   XOR2_X1 U412 (.A(RF_OUT2[14]),
	.B(RF_OUT1[14]),
	.Z(n303));
   XOR2_X1 U413 (.A(RF_OUT2[13]),
	.B(RF_OUT1[13]),
	.Z(n302));
   XOR2_X1 U414 (.A(RF_OUT2[12]),
	.B(RF_OUT1[12]),
	.Z(n301));
   XOR2_X1 U415 (.A(RF_OUT2[11]),
	.B(RF_OUT1[11]),
	.Z(n316));
   XOR2_X1 U416 (.A(RF_OUT2[10]),
	.B(RF_OUT1[10]),
	.Z(n315));
   XOR2_X1 U417 (.A(RF_OUT2[9]),
	.B(RF_OUT1[9]),
	.Z(n314));
   XOR2_X1 U418 (.A(RF_OUT2[8]),
	.B(RF_OUT1[8]),
	.Z(n313));
   XOR2_X1 U419 (.A(RF_OUT2[7]),
	.B(RF_OUT1[7]),
	.Z(n328));
   XOR2_X1 U420 (.A(RF_OUT2[6]),
	.B(RF_OUT1[6]),
	.Z(n327));
   XOR2_X1 U421 (.A(RF_OUT2[5]),
	.B(RF_OUT1[5]),
	.Z(n326));
   XOR2_X1 U422 (.A(RF_OUT2[4]),
	.B(RF_OUT1[4]),
	.Z(n325));
   XOR2_X1 U423 (.A(RF_OUT2[3]),
	.B(RF_OUT1[3]),
	.Z(n340));
   XOR2_X1 U424 (.A(RF_OUT2[2]),
	.B(RF_OUT1[2]),
	.Z(n339));
   XOR2_X1 U425 (.A(RF_OUT2[1]),
	.B(RF_OUT1[1]),
	.Z(n338));
   XOR2_X1 U426 (.A(RF_OUT2[0]),
	.B(RF_OUT1[0]),
	.Z(n337));
   NAND3_X1 U428 (.A1(n384),
	.A2(n385),
	.A3(MUX_IMM_SEL[1]),
	.ZN(n356));
   register_file_NBITS32 rf (.CLK(clk),
	.RESET(rst),
	.ENABLE(en),
	.RD1(RF_RD1),
	.RD2(RF_RD2),
	.WR(RF_WR),
	.ADD_WR(ADD_WR),
	.ADD_RD1(RS1),
	.ADD_RD2(RS2),
	.DATAIN(DATAIN),
	.OUT1(RF_OUT1_m),
	.OUT2(RF_OUT2_m));
   decode_unit_DW01_add_0 add_123 (.A(PC_OUT),
	.B(IMM),
	.CI(1'b0),
	.SUM(JMP_ADDR));
   DFF_X1 currIR_reg_3_ (.D(n92),
	.CK(clk),
	.Q(OPCODE[3]));
   DFF_X1 currIR_reg_1_ (.D(n94),
	.CK(clk),
	.Q(OPCODE[1]));
   DFF_X1 currIR_reg_0_ (.D(n95),
	.CK(clk),
	.Q(OPCODE[0]),
	.QN(n6));
   NOR2_X1 U3 (.A1(n349),
	.A2(n51),
	.ZN(IMM[5]));
   INV_X1 U5 (.A(n8),
	.ZN(n357));
   OAI21_X1 U6 (.A(n352),
	.B1(n59),
	.B2(n383),
	.ZN(IMM[21]));
   OAI21_X1 U7 (.A(n352),
	.B1(n53),
	.B2(n383),
	.ZN(IMM[24]));
   OAI21_X1 U8 (.A(n352),
	.B1(n51),
	.B2(n383),
	.ZN(IMM[25]));
   OAI21_X1 U9 (.A(n352),
	.B1(n43),
	.B2(n383),
	.ZN(IMM[29]));
   OAI21_X1 U10 (.A(n352),
	.B1(n41),
	.B2(n383),
	.ZN(IMM[30]));
   OAI22_X1 U12 (.A1(n350),
	.A2(n59),
	.B1(n351),
	.B2(n85),
	.ZN(IMM[1]));
   OR3_X1 U13 (.A1(MUX_IMM_SEL[1]),
	.A2(MUX_IMM_SEL[2]),
	.A3(MUX_IMM_SEL[0]),
	.ZN(n4));
   INV_X1 U15 (.A(n6),
	.ZN(n7));
   OR3_X1 U16 (.A1(MUX_IMM_SEL[1]),
	.A2(MUX_IMM_SEL[2]),
	.A3(n384),
	.ZN(n9));
   AND3_X1 U17 (.A1(MUX_IMM_SEL[0]),
	.A2(n385),
	.A3(MUX_IMM_SEL[1]),
	.ZN(n8));
   INV_X1 U18 (.A(n9),
	.ZN(n359));
   NOR2_X1 U19 (.A1(n354),
	.A2(n8),
	.ZN(n349));
   NOR2_X1 U20 (.A1(n353),
	.A2(n8),
	.ZN(n350));
   INV_X1 U21 (.A(n349),
	.ZN(n383));
   NAND4_X1 U28 (.A1(n239),
	.A2(n240),
	.A3(n241),
	.A4(n242),
	.ZN(n238));
   NOR4_X1 U29 (.A1(n285),
	.A2(n286),
	.A3(n287),
	.A4(n288),
	.ZN(n239));
   NOR4_X1 U30 (.A1(n261),
	.A2(n262),
	.A3(n263),
	.A4(n264),
	.ZN(n241));
   NOR4_X1 U31 (.A1(n243),
	.A2(n244),
	.A3(n245),
	.A4(n246),
	.ZN(n242));
   NOR3_X1 U32 (.A1(MUX_IMM_SEL[1]),
	.A2(MUX_IMM_SEL[2]),
	.A3(MUX_IMM_SEL[0]),
	.ZN(n353));
   INV_X1 U33 (.A(MUX_IMM_SEL[2]),
	.ZN(n385));
   INV_X1 U34 (.A(MUX_IMM_SEL[0]),
	.ZN(n384));
   NOR4_X1 U37 (.A1(n301),
	.A2(n302),
	.A3(n303),
	.A4(n304),
	.ZN(n300));
   NOR4_X1 U38 (.A1(n313),
	.A2(n314),
	.A3(n315),
	.A4(n316),
	.ZN(n299));
   NOR4_X1 U39 (.A1(n273),
	.A2(n274),
	.A3(n275),
	.A4(n276),
	.ZN(n240));
   NOR4_X1 U40 (.A1(n325),
	.A2(n326),
	.A3(n327),
	.A4(n328),
	.ZN(n298));
   NOR4_X1 U41 (.A1(n337),
	.A2(n338),
	.A3(n339),
	.A4(n340),
	.ZN(n297));
   NAND2_X2 U50 (.A1(n247),
	.A2(n10),
	.ZN(n248));
   NAND2_X2 U51 (.A1(n251),
	.A2(n11),
	.ZN(n252));
   OAI221_X1 U52 (.A(n329),
	.B1(n375),
	.B2(n247),
	.C1(n122),
	.C2(n248),
	.ZN(RF_OUT1[7]));
   NAND2_X1 U53 (.A1(RF_OUT1_m[7]),
	.A2(FE_DBTN2_n10),
	.ZN(n329));
   OAI221_X1 U54 (.A(n331),
	.B1(n376),
	.B2(n247),
	.C1(n123),
	.C2(n248),
	.ZN(RF_OUT1[6]));
   NAND2_X1 U55 (.A1(RF_OUT1_m[6]),
	.A2(FE_DBTN2_n10),
	.ZN(n331));
   OAI221_X1 U56 (.A(n333),
	.B1(n377),
	.B2(n247),
	.C1(n124),
	.C2(n248),
	.ZN(RF_OUT1[5]));
   NAND2_X1 U57 (.A1(RF_OUT1_m[5]),
	.A2(FE_DBTN2_n10),
	.ZN(n333));
   OAI221_X1 U58 (.A(n335),
	.B1(n378),
	.B2(n247),
	.C1(n125),
	.C2(n248),
	.ZN(RF_OUT1[4]));
   NAND2_X1 U59 (.A1(RF_OUT1_m[4]),
	.A2(FE_DBTN2_n10),
	.ZN(n335));
   OAI221_X1 U60 (.A(n341),
	.B1(n379),
	.B2(n247),
	.C1(n126),
	.C2(n248),
	.ZN(RF_OUT1[3]));
   NAND2_X1 U61 (.A1(RF_OUT1_m[3]),
	.A2(FE_DBTN2_n10),
	.ZN(n341));
   OAI221_X1 U62 (.A(n343),
	.B1(n380),
	.B2(n247),
	.C1(n127),
	.C2(n248),
	.ZN(RF_OUT1[2]));
   NAND2_X1 U63 (.A1(RF_OUT1_m[2]),
	.A2(FE_DBTN2_n10),
	.ZN(n343));
   OAI221_X1 U64 (.A(n345),
	.B1(n381),
	.B2(n247),
	.C1(n128),
	.C2(n248),
	.ZN(RF_OUT1[1]));
   NAND2_X1 U65 (.A1(RF_OUT1_m[1]),
	.A2(FE_DBTN2_n10),
	.ZN(n345));
   OAI221_X1 U66 (.A(n347),
	.B1(n382),
	.B2(n247),
	.C1(n129),
	.C2(n248),
	.ZN(RF_OUT1[0]));
   NAND2_X1 U67 (.A1(RF_OUT1_m[0]),
	.A2(FE_DBTN2_n10),
	.ZN(n347));
   OAI221_X1 U68 (.A(n277),
	.B1(n254),
	.B2(n247),
	.C1(n106),
	.C2(n248),
	.ZN(RF_OUT1[23]));
   NAND2_X1 U69 (.A1(RF_OUT1_m[23]),
	.A2(FE_DBTN2_n10),
	.ZN(n277));
   OAI221_X1 U70 (.A(n279),
	.B1(n360),
	.B2(n247),
	.C1(n107),
	.C2(n248),
	.ZN(RF_OUT1[22]));
   NAND2_X1 U71 (.A1(RF_OUT1_m[22]),
	.A2(FE_DBTN2_n10),
	.ZN(n279));
   OAI221_X1 U72 (.A(n281),
	.B1(n361),
	.B2(n247),
	.C1(n108),
	.C2(n248),
	.ZN(RF_OUT1[21]));
   NAND2_X1 U73 (.A1(RF_OUT1_m[21]),
	.A2(FE_DBTN2_n10),
	.ZN(n281));
   OAI221_X1 U74 (.A(n283),
	.B1(n362),
	.B2(n247),
	.C1(n109),
	.C2(n248),
	.ZN(RF_OUT1[20]));
   NAND2_X1 U75 (.A1(RF_OUT1_m[20]),
	.A2(FE_DBTN2_n10),
	.ZN(n283));
   OAI221_X1 U76 (.A(n249),
	.B1(n162),
	.B2(n247),
	.C1(n98),
	.C2(n248),
	.ZN(RF_OUT1[31]));
   NAND2_X1 U77 (.A1(RF_OUT1_m[31]),
	.A2(FE_DBTN2_n10),
	.ZN(n249));
   OAI221_X1 U78 (.A(n255),
	.B1(n163),
	.B2(n247),
	.C1(n99),
	.C2(n248),
	.ZN(RF_OUT1[30]));
   NAND2_X1 U79 (.A1(RF_OUT1_m[30]),
	.A2(FE_DBTN2_n10),
	.ZN(n255));
   OAI221_X1 U80 (.A(n257),
	.B1(n164),
	.B2(n247),
	.C1(n100),
	.C2(n248),
	.ZN(RF_OUT1[29]));
   NAND2_X1 U81 (.A1(RF_OUT1_m[29]),
	.A2(FE_DBTN2_n10),
	.ZN(n257));
   OAI221_X1 U82 (.A(n259),
	.B1(n165),
	.B2(n247),
	.C1(n101),
	.C2(n248),
	.ZN(RF_OUT1[28]));
   NAND2_X1 U83 (.A1(RF_OUT1_m[28]),
	.A2(FE_DBTN2_n10),
	.ZN(n259));
   OAI221_X1 U84 (.A(n265),
	.B1(n166),
	.B2(n247),
	.C1(n102),
	.C2(n248),
	.ZN(RF_OUT1[27]));
   NAND2_X1 U85 (.A1(RF_OUT1_m[27]),
	.A2(FE_DBTN2_n10),
	.ZN(n265));
   OAI221_X1 U86 (.A(n267),
	.B1(n167),
	.B2(n247),
	.C1(n103),
	.C2(n248),
	.ZN(RF_OUT1[26]));
   NAND2_X1 U87 (.A1(RF_OUT1_m[26]),
	.A2(FE_DBTN2_n10),
	.ZN(n267));
   OAI221_X1 U88 (.A(n269),
	.B1(n168),
	.B2(n247),
	.C1(n104),
	.C2(n248),
	.ZN(RF_OUT1[25]));
   NAND2_X1 U89 (.A1(RF_OUT1_m[25]),
	.A2(FE_DBTN2_n10),
	.ZN(n269));
   OAI221_X1 U90 (.A(n271),
	.B1(n250),
	.B2(n247),
	.C1(n105),
	.C2(n248),
	.ZN(RF_OUT1[24]));
   NAND2_X1 U91 (.A1(RF_OUT1_m[24]),
	.A2(FE_DBTN2_n10),
	.ZN(n271));
   OAI221_X1 U92 (.A(n289),
	.B1(n363),
	.B2(n247),
	.C1(n110),
	.C2(n248),
	.ZN(RF_OUT1[19]));
   NAND2_X1 U93 (.A1(RF_OUT1_m[19]),
	.A2(FE_DBTN2_n10),
	.ZN(n289));
   OAI221_X1 U94 (.A(n291),
	.B1(n364),
	.B2(n247),
	.C1(n111),
	.C2(n248),
	.ZN(RF_OUT1[18]));
   NAND2_X1 U95 (.A1(RF_OUT1_m[18]),
	.A2(FE_DBTN2_n10),
	.ZN(n291));
   OAI221_X1 U96 (.A(n293),
	.B1(n365),
	.B2(n247),
	.C1(n112),
	.C2(n248),
	.ZN(RF_OUT1[17]));
   NAND2_X1 U97 (.A1(RF_OUT1_m[17]),
	.A2(FE_DBTN2_n10),
	.ZN(n293));
   OAI221_X1 U98 (.A(n295),
	.B1(n366),
	.B2(n247),
	.C1(n113),
	.C2(n248),
	.ZN(RF_OUT1[16]));
   NAND2_X1 U99 (.A1(RF_OUT1_m[16]),
	.A2(FE_DBTN2_n10),
	.ZN(n295));
   OAI221_X1 U100 (.A(n305),
	.B1(n367),
	.B2(n247),
	.C1(n114),
	.C2(n248),
	.ZN(RF_OUT1[15]));
   NAND2_X1 U101 (.A1(RF_OUT1_m[15]),
	.A2(FE_DBTN2_n10),
	.ZN(n305));
   OAI221_X1 U102 (.A(n307),
	.B1(n368),
	.B2(n247),
	.C1(n115),
	.C2(n248),
	.ZN(RF_OUT1[14]));
   NAND2_X1 U103 (.A1(RF_OUT1_m[14]),
	.A2(FE_DBTN2_n10),
	.ZN(n307));
   OAI221_X1 U104 (.A(n309),
	.B1(n369),
	.B2(n247),
	.C1(n116),
	.C2(n248),
	.ZN(RF_OUT1[13]));
   NAND2_X1 U105 (.A1(RF_OUT1_m[13]),
	.A2(FE_DBTN2_n10),
	.ZN(n309));
   OAI221_X1 U106 (.A(n311),
	.B1(n370),
	.B2(n247),
	.C1(n117),
	.C2(n248),
	.ZN(RF_OUT1[12]));
   NAND2_X1 U107 (.A1(RF_OUT1_m[12]),
	.A2(FE_DBTN2_n10),
	.ZN(n311));
   OAI221_X1 U108 (.A(n317),
	.B1(n371),
	.B2(n247),
	.C1(n118),
	.C2(n248),
	.ZN(RF_OUT1[11]));
   NAND2_X1 U109 (.A1(RF_OUT1_m[11]),
	.A2(FE_DBTN2_n10),
	.ZN(n317));
   OAI221_X1 U110 (.A(n319),
	.B1(n372),
	.B2(n247),
	.C1(n119),
	.C2(n248),
	.ZN(RF_OUT1[10]));
   NAND2_X1 U111 (.A1(RF_OUT1_m[10]),
	.A2(FE_DBTN2_n10),
	.ZN(n319));
   OAI221_X1 U112 (.A(n321),
	.B1(n373),
	.B2(n247),
	.C1(n120),
	.C2(n248),
	.ZN(RF_OUT1[9]));
   NAND2_X1 U113 (.A1(RF_OUT1_m[9]),
	.A2(FE_DBTN2_n10),
	.ZN(n321));
   OAI221_X1 U114 (.A(n323),
	.B1(n374),
	.B2(n247),
	.C1(n121),
	.C2(n248),
	.ZN(RF_OUT1[8]));
   NAND2_X1 U115 (.A1(RF_OUT1_m[8]),
	.A2(FE_DBTN2_n10),
	.ZN(n323));
   OAI221_X1 U116 (.A(n278),
	.B1(n251),
	.B2(n254),
	.C1(n252),
	.C2(n106),
	.ZN(RF_OUT2[23]));
   NAND2_X1 U117 (.A1(RF_OUT2_m[23]),
	.A2(FE_DBTN1_n11),
	.ZN(n278));
   OAI221_X1 U118 (.A(n280),
	.B1(n251),
	.B2(n360),
	.C1(n252),
	.C2(n107),
	.ZN(RF_OUT2[22]));
   NAND2_X1 U119 (.A1(RF_OUT2_m[22]),
	.A2(FE_DBTN1_n11),
	.ZN(n280));
   OAI221_X1 U120 (.A(n282),
	.B1(n251),
	.B2(n361),
	.C1(n252),
	.C2(n108),
	.ZN(RF_OUT2[21]));
   NAND2_X1 U121 (.A1(RF_OUT2_m[21]),
	.A2(FE_DBTN1_n11),
	.ZN(n282));
   OAI221_X1 U122 (.A(n284),
	.B1(n251),
	.B2(n362),
	.C1(n252),
	.C2(n109),
	.ZN(RF_OUT2[20]));
   NAND2_X1 U123 (.A1(RF_OUT2_m[20]),
	.A2(FE_DBTN1_n11),
	.ZN(n284));
   OAI221_X1 U124 (.A(n253),
	.B1(n251),
	.B2(n162),
	.C1(n252),
	.C2(n98),
	.ZN(RF_OUT2[31]));
   NAND2_X1 U125 (.A1(RF_OUT2_m[31]),
	.A2(FE_DBTN1_n11),
	.ZN(n253));
   OAI221_X1 U126 (.A(n256),
	.B1(n251),
	.B2(n163),
	.C1(n252),
	.C2(n99),
	.ZN(RF_OUT2[30]));
   NAND2_X1 U127 (.A1(RF_OUT2_m[30]),
	.A2(FE_DBTN1_n11),
	.ZN(n256));
   OAI221_X1 U128 (.A(n258),
	.B1(n251),
	.B2(n164),
	.C1(n252),
	.C2(n100),
	.ZN(RF_OUT2[29]));
   NAND2_X1 U129 (.A1(RF_OUT2_m[29]),
	.A2(FE_DBTN1_n11),
	.ZN(n258));
   OAI221_X1 U130 (.A(n260),
	.B1(n251),
	.B2(n165),
	.C1(n252),
	.C2(n101),
	.ZN(RF_OUT2[28]));
   NAND2_X1 U131 (.A1(RF_OUT2_m[28]),
	.A2(FE_DBTN1_n11),
	.ZN(n260));
   OAI221_X1 U132 (.A(n266),
	.B1(n251),
	.B2(n166),
	.C1(n252),
	.C2(n102),
	.ZN(RF_OUT2[27]));
   NAND2_X1 U133 (.A1(RF_OUT2_m[27]),
	.A2(FE_DBTN1_n11),
	.ZN(n266));
   OAI221_X1 U134 (.A(n268),
	.B1(n251),
	.B2(n167),
	.C1(n252),
	.C2(n103),
	.ZN(RF_OUT2[26]));
   NAND2_X1 U135 (.A1(RF_OUT2_m[26]),
	.A2(FE_DBTN1_n11),
	.ZN(n268));
   OAI221_X1 U136 (.A(n270),
	.B1(n251),
	.B2(n168),
	.C1(n252),
	.C2(n104),
	.ZN(RF_OUT2[25]));
   NAND2_X1 U137 (.A1(RF_OUT2_m[25]),
	.A2(FE_DBTN1_n11),
	.ZN(n270));
   OAI221_X1 U138 (.A(n272),
	.B1(n251),
	.B2(n250),
	.C1(n252),
	.C2(n105),
	.ZN(RF_OUT2[24]));
   NAND2_X1 U139 (.A1(RF_OUT2_m[24]),
	.A2(FE_DBTN1_n11),
	.ZN(n272));
   OAI221_X1 U140 (.A(n290),
	.B1(n251),
	.B2(n363),
	.C1(n252),
	.C2(n110),
	.ZN(RF_OUT2[19]));
   NAND2_X1 U141 (.A1(RF_OUT2_m[19]),
	.A2(FE_DBTN1_n11),
	.ZN(n290));
   OAI221_X1 U142 (.A(n292),
	.B1(n251),
	.B2(n364),
	.C1(n252),
	.C2(n111),
	.ZN(RF_OUT2[18]));
   NAND2_X1 U143 (.A1(RF_OUT2_m[18]),
	.A2(FE_DBTN1_n11),
	.ZN(n292));
   OAI221_X1 U144 (.A(n294),
	.B1(n251),
	.B2(n365),
	.C1(n252),
	.C2(n112),
	.ZN(RF_OUT2[17]));
   NAND2_X1 U145 (.A1(RF_OUT2_m[17]),
	.A2(FE_DBTN1_n11),
	.ZN(n294));
   OAI221_X1 U146 (.A(n296),
	.B1(n251),
	.B2(n366),
	.C1(n252),
	.C2(n113),
	.ZN(RF_OUT2[16]));
   NAND2_X1 U147 (.A1(RF_OUT2_m[16]),
	.A2(FE_DBTN1_n11),
	.ZN(n296));
   OAI221_X1 U148 (.A(n306),
	.B1(n251),
	.B2(n367),
	.C1(n252),
	.C2(n114),
	.ZN(RF_OUT2[15]));
   NAND2_X1 U149 (.A1(RF_OUT2_m[15]),
	.A2(FE_DBTN1_n11),
	.ZN(n306));
   OAI221_X1 U150 (.A(n308),
	.B1(n251),
	.B2(n368),
	.C1(n252),
	.C2(n115),
	.ZN(RF_OUT2[14]));
   NAND2_X1 U151 (.A1(RF_OUT2_m[14]),
	.A2(FE_DBTN1_n11),
	.ZN(n308));
   OAI221_X1 U152 (.A(n310),
	.B1(n251),
	.B2(n369),
	.C1(n252),
	.C2(n116),
	.ZN(RF_OUT2[13]));
   NAND2_X1 U153 (.A1(RF_OUT2_m[13]),
	.A2(FE_DBTN1_n11),
	.ZN(n310));
   OAI221_X1 U154 (.A(n312),
	.B1(n251),
	.B2(n370),
	.C1(n252),
	.C2(n117),
	.ZN(RF_OUT2[12]));
   NAND2_X1 U155 (.A1(RF_OUT2_m[12]),
	.A2(FE_DBTN1_n11),
	.ZN(n312));
   OAI221_X1 U156 (.A(n318),
	.B1(n251),
	.B2(n371),
	.C1(n252),
	.C2(n118),
	.ZN(RF_OUT2[11]));
   NAND2_X1 U157 (.A1(RF_OUT2_m[11]),
	.A2(FE_DBTN1_n11),
	.ZN(n318));
   OAI221_X1 U158 (.A(n320),
	.B1(n251),
	.B2(n372),
	.C1(n252),
	.C2(n119),
	.ZN(RF_OUT2[10]));
   NAND2_X1 U159 (.A1(RF_OUT2_m[10]),
	.A2(FE_DBTN1_n11),
	.ZN(n320));
   OAI221_X1 U160 (.A(n322),
	.B1(n251),
	.B2(n373),
	.C1(n252),
	.C2(n120),
	.ZN(RF_OUT2[9]));
   NAND2_X1 U161 (.A1(RF_OUT2_m[9]),
	.A2(FE_DBTN1_n11),
	.ZN(n322));
   OAI221_X1 U162 (.A(n324),
	.B1(n251),
	.B2(n374),
	.C1(n252),
	.C2(n121),
	.ZN(RF_OUT2[8]));
   NAND2_X1 U163 (.A1(RF_OUT2_m[8]),
	.A2(FE_DBTN1_n11),
	.ZN(n324));
   OAI221_X1 U164 (.A(n330),
	.B1(n251),
	.B2(n375),
	.C1(n252),
	.C2(n122),
	.ZN(RF_OUT2[7]));
   NAND2_X1 U165 (.A1(RF_OUT2_m[7]),
	.A2(FE_DBTN1_n11),
	.ZN(n330));
   OAI221_X1 U166 (.A(n332),
	.B1(n251),
	.B2(n376),
	.C1(n252),
	.C2(n123),
	.ZN(RF_OUT2[6]));
   NAND2_X1 U167 (.A1(RF_OUT2_m[6]),
	.A2(FE_DBTN1_n11),
	.ZN(n332));
   OAI221_X1 U168 (.A(n334),
	.B1(n251),
	.B2(n377),
	.C1(n252),
	.C2(n124),
	.ZN(RF_OUT2[5]));
   NAND2_X1 U169 (.A1(RF_OUT2_m[5]),
	.A2(FE_DBTN1_n11),
	.ZN(n334));
   OAI221_X1 U170 (.A(n336),
	.B1(n251),
	.B2(n378),
	.C1(n252),
	.C2(n125),
	.ZN(RF_OUT2[4]));
   NAND2_X1 U171 (.A1(RF_OUT2_m[4]),
	.A2(FE_DBTN1_n11),
	.ZN(n336));
   OAI221_X1 U172 (.A(n342),
	.B1(n251),
	.B2(n379),
	.C1(n252),
	.C2(n126),
	.ZN(RF_OUT2[3]));
   NAND2_X1 U173 (.A1(RF_OUT2_m[3]),
	.A2(FE_DBTN1_n11),
	.ZN(n342));
   OAI221_X1 U174 (.A(n344),
	.B1(n251),
	.B2(n380),
	.C1(n252),
	.C2(n127),
	.ZN(RF_OUT2[2]));
   NAND2_X1 U175 (.A1(RF_OUT2_m[2]),
	.A2(FE_DBTN1_n11),
	.ZN(n344));
   OAI221_X1 U176 (.A(n346),
	.B1(n251),
	.B2(n381),
	.C1(n252),
	.C2(n128),
	.ZN(RF_OUT2[1]));
   NAND2_X1 U177 (.A1(RF_OUT2_m[1]),
	.A2(FE_DBTN1_n11),
	.ZN(n346));
   OAI221_X1 U178 (.A(n348),
	.B1(n251),
	.B2(n382),
	.C1(n252),
	.C2(n129),
	.ZN(RF_OUT2[0]));
   NAND2_X1 U179 (.A1(RF_OUT2_m[0]),
	.A2(FE_DBTN1_n11),
	.ZN(n348));
   NOR2_X1 U185 (.A1(n237),
	.A2(n238),
	.ZN(EQU_FLAG));
   NAND4_X1 U186 (.A1(n297),
	.A2(n298),
	.A3(n299),
	.A4(n300),
	.ZN(n237));
   OR2_X1 U187 (.A1(RF_OUT1_SEL[1]),
	.A2(RF_OUT1_SEL[0]),
	.ZN(n10));
   OR2_X1 U188 (.A1(RF_OUT2_SEL[1]),
	.A2(RF_OUT2_SEL[0]),
	.ZN(n11));
   NAND2_X2 U189 (.A1(RF_OUT2_SEL[0]),
	.A2(n96),
	.ZN(n251));
   INV_X1 U190 (.A(RF_OUT2_SEL[1]),
	.ZN(n96));
   NAND2_X2 U192 (.A1(RF_OUT1_SEL[0]),
	.A2(n97),
	.ZN(n247));
   INV_X1 U193 (.A(RF_OUT1_SEL[1]),
	.ZN(n97));
   INV_X1 U194 (.A(DATAIN[31]),
	.ZN(n98));
   INV_X1 U195 (.A(DATAIN[23]),
	.ZN(n106));
   INV_X1 U196 (.A(DATAIN[22]),
	.ZN(n107));
   INV_X1 U197 (.A(DATAIN[21]),
	.ZN(n108));
   INV_X1 U198 (.A(DATAIN[20]),
	.ZN(n109));
   INV_X1 U199 (.A(DATAIN[30]),
	.ZN(n99));
   INV_X1 U200 (.A(DATAIN[29]),
	.ZN(n100));
   INV_X1 U201 (.A(DATAIN[28]),
	.ZN(n101));
   INV_X1 U202 (.A(DATAIN[27]),
	.ZN(n102));
   INV_X1 U203 (.A(DATAIN[26]),
	.ZN(n103));
   INV_X1 U204 (.A(DATAIN[25]),
	.ZN(n104));
   INV_X1 U205 (.A(DATAIN[24]),
	.ZN(n105));
   INV_X1 U206 (.A(DATAIN[2]),
	.ZN(n127));
   INV_X1 U207 (.A(DATAIN[9]),
	.ZN(n120));
   INV_X1 U208 (.A(DATAIN[8]),
	.ZN(n121));
   INV_X1 U209 (.A(DATAIN[7]),
	.ZN(n122));
   INV_X1 U210 (.A(DATAIN[6]),
	.ZN(n123));
   INV_X1 U211 (.A(DATAIN[5]),
	.ZN(n124));
   INV_X1 U212 (.A(DATAIN[4]),
	.ZN(n125));
   INV_X1 U213 (.A(DATAIN[3]),
	.ZN(n126));
   INV_X1 U214 (.A(DATAIN[19]),
	.ZN(n110));
   INV_X1 U215 (.A(DATAIN[18]),
	.ZN(n111));
   INV_X1 U216 (.A(DATAIN[17]),
	.ZN(n112));
   INV_X1 U217 (.A(DATAIN[16]),
	.ZN(n113));
   INV_X1 U218 (.A(DATAIN[15]),
	.ZN(n114));
   INV_X1 U219 (.A(DATAIN[14]),
	.ZN(n115));
   INV_X1 U220 (.A(DATAIN[13]),
	.ZN(n116));
   INV_X1 U221 (.A(DATAIN[12]),
	.ZN(n117));
   INV_X1 U222 (.A(DATAIN[11]),
	.ZN(n118));
   INV_X1 U223 (.A(DATAIN[10]),
	.ZN(n119));
   INV_X1 U224 (.A(DATAIN[1]),
	.ZN(n128));
   INV_X1 U225 (.A(DATAIN[0]),
	.ZN(n129));
   NAND2_X1 U232 (.A1(IMM[31]),
	.A2(n383),
	.ZN(n352));
   OAI22_X1 U233 (.A1(n61),
	.A2(n4),
	.B1(n87),
	.B2(n9),
	.ZN(IMM[0]));
   OAI221_X1 U234 (.A(n358),
	.B1(n87),
	.B2(n356),
	.C1(n61),
	.C2(n357),
	.ZN(IMM[11]));
   OAI21_X1 U235 (.A(IMM[31]),
	.B1(n353),
	.B2(n359),
	.ZN(n358));
   OAI22_X1 U237 (.A1(n350),
	.A2(n53),
	.B1(n351),
	.B2(n79),
	.ZN(IMM[4]));
   OAI22_X1 U238 (.A1(n350),
	.A2(n55),
	.B1(n351),
	.B2(n81),
	.ZN(IMM[3]));
   OAI22_X1 U239 (.A1(n350),
	.A2(n57),
	.B1(n351),
	.B2(n83),
	.ZN(IMM[2]));
   NAND2_X1 U240 (.A1(IMM[31]),
	.A2(n354),
	.ZN(n355));
   OAI21_X1 U241 (.A(n355),
	.B1(n75),
	.B2(n354),
	.ZN(IMM[13]));
   OAI21_X1 U242 (.A(n355),
	.B1(n77),
	.B2(n354),
	.ZN(IMM[12]));
   OAI21_X1 U243 (.A(n355),
	.B1(n73),
	.B2(n354),
	.ZN(IMM[14]));
   OAI21_X1 U244 (.A(n355),
	.B1(n71),
	.B2(n354),
	.ZN(IMM[15]));
   OAI21_X1 U245 (.A(n355),
	.B1(n69),
	.B2(n354),
	.ZN(IMM[16]));
   OAI21_X1 U246 (.A(n355),
	.B1(n67),
	.B2(n354),
	.ZN(IMM[17]));
   OAI21_X1 U247 (.A(n355),
	.B1(n65),
	.B2(n354),
	.ZN(IMM[18]));
   OAI21_X1 U248 (.A(n355),
	.B1(n63),
	.B2(n354),
	.ZN(IMM[19]));
   OAI21_X1 U249 (.A(n352),
	.B1(n61),
	.B2(n383),
	.ZN(IMM[20]));
   OAI21_X1 U250 (.A(n352),
	.B1(n57),
	.B2(n383),
	.ZN(IMM[22]));
   OAI21_X1 U251 (.A(n352),
	.B1(n55),
	.B2(n383),
	.ZN(IMM[23]));
   NOR2_X1 U254 (.A1(n349),
	.A2(n45),
	.ZN(IMM[8]));
   NOR2_X1 U255 (.A1(n349),
	.A2(n43),
	.ZN(IMM[9]));
   NOR2_X1 U256 (.A1(n349),
	.A2(n47),
	.ZN(IMM[7]));
   NOR2_X1 U257 (.A1(n349),
	.A2(n49),
	.ZN(IMM[6]));
   NOR2_X1 U258 (.A1(n349),
	.A2(n41),
	.ZN(IMM[10]));
   NOR3_X1 U259 (.A1(IF_FLUSH),
	.A2(rst),
	.A3(FE_OFN29_n171),
	.ZN(n170));
   NOR3_X1 U260 (.A1(en),
	.A2(rst),
	.A3(IF_FLUSH),
	.ZN(n171));
   OAI21_X1 U261 (.A(n352),
	.B1(n49),
	.B2(n383),
	.ZN(IMM[26]));
   OAI21_X1 U262 (.A(n352),
	.B1(n47),
	.B2(n383),
	.ZN(IMM[27]));
   OAI21_X1 U263 (.A(n352),
	.B1(n45),
	.B2(n383),
	.ZN(IMM[28]));
   INV_X1 U264 (.A(n172),
	.ZN(n94));
   AOI22_X1 U265 (.A1(IR_IN[1]),
	.A2(FE_OFN92_n170),
	.B1(OPCODE[1]),
	.B2(FE_OFN29_n171),
	.ZN(n172));
   INV_X1 U266 (.A(n184),
	.ZN(n76));
   AOI22_X1 U267 (.A1(FE_OFN29_n171),
	.A2(FUNC3[1]),
	.B1(FE_OFN92_n170),
	.B2(IR_IN[13]),
	.ZN(n184));
   INV_X1 U268 (.A(n185),
	.ZN(n74));
   AOI22_X1 U269 (.A1(FE_OFN29_n171),
	.A2(FUNC3[2]),
	.B1(FE_OFN92_n170),
	.B2(IR_IN[14]),
	.ZN(n185));
   INV_X1 U270 (.A(n196),
	.ZN(n52));
   AOI22_X1 U271 (.A1(FE_OFN29_n171),
	.A2(currIR[25]),
	.B1(FE_OFN92_n170),
	.B2(IR_IN[25]),
	.ZN(n196));
   INV_X1 U272 (.A(n197),
	.ZN(n50));
   AOI22_X1 U273 (.A1(FE_OFN29_n171),
	.A2(currIR[26]),
	.B1(FE_OFN92_n170),
	.B2(IR_IN[26]),
	.ZN(n197));
   INV_X1 U274 (.A(n198),
	.ZN(n48));
   AOI22_X1 U275 (.A1(FE_OFN29_n171),
	.A2(currIR[27]),
	.B1(FE_OFN92_n170),
	.B2(IR_IN[27]),
	.ZN(n198));
   INV_X1 U276 (.A(n199),
	.ZN(n46));
   AOI22_X1 U277 (.A1(FE_OFN29_n171),
	.A2(currIR[28]),
	.B1(FE_OFN92_n170),
	.B2(IR_IN[28]),
	.ZN(n199));
   INV_X1 U278 (.A(n200),
	.ZN(n44));
   AOI22_X1 U279 (.A1(FE_OFN29_n171),
	.A2(currIR[29]),
	.B1(FE_OFN92_n170),
	.B2(IR_IN[29]),
	.ZN(n200));
   INV_X1 U280 (.A(n201),
	.ZN(n42));
   AOI22_X1 U281 (.A1(FE_OFN29_n171),
	.A2(currIR[30]),
	.B1(FE_OFN92_n170),
	.B2(IR_IN[30]),
	.ZN(n201));
   INV_X1 U282 (.A(EXE_MEM_IN[2]),
	.ZN(n380));
   INV_X1 U283 (.A(EXE_MEM_IN[23]),
	.ZN(n254));
   INV_X1 U284 (.A(EXE_MEM_IN[22]),
	.ZN(n360));
   INV_X1 U285 (.A(EXE_MEM_IN[21]),
	.ZN(n361));
   INV_X1 U286 (.A(EXE_MEM_IN[30]),
	.ZN(n163));
   INV_X1 U287 (.A(EXE_MEM_IN[29]),
	.ZN(n164));
   INV_X1 U288 (.A(EXE_MEM_IN[27]),
	.ZN(n166));
   INV_X1 U289 (.A(EXE_MEM_IN[26]),
	.ZN(n167));
   INV_X1 U290 (.A(EXE_MEM_IN[25]),
	.ZN(n168));
   INV_X1 U291 (.A(EXE_MEM_IN[19]),
	.ZN(n363));
   INV_X1 U292 (.A(EXE_MEM_IN[18]),
	.ZN(n364));
   INV_X1 U293 (.A(EXE_MEM_IN[15]),
	.ZN(n367));
   INV_X1 U294 (.A(EXE_MEM_IN[14]),
	.ZN(n368));
   INV_X1 U295 (.A(EXE_MEM_IN[11]),
	.ZN(n371));
   INV_X1 U296 (.A(EXE_MEM_IN[10]),
	.ZN(n372));
   INV_X1 U297 (.A(EXE_MEM_IN[7]),
	.ZN(n375));
   INV_X1 U298 (.A(EXE_MEM_IN[6]),
	.ZN(n376));
   INV_X1 U299 (.A(EXE_MEM_IN[3]),
	.ZN(n379));
   INV_X1 U300 (.A(EXE_MEM_IN[31]),
	.ZN(n162));
   INV_X1 U301 (.A(n173),
	.ZN(n93));
   AOI22_X1 U302 (.A1(IR_IN[2]),
	.A2(FE_OFN92_n170),
	.B1(OPCODE[2]),
	.B2(FE_OFN29_n171),
	.ZN(n173));
   INV_X1 U303 (.A(n169),
	.ZN(n95));
   INV_X1 U304 (.A(n188),
	.ZN(n68));
   AOI22_X1 U305 (.A1(FE_OFN29_n171),
	.A2(RS1[2]),
	.B1(FE_OFN92_n170),
	.B2(IR_IN[17]),
	.ZN(n188));
   INV_X1 U306 (.A(n193),
	.ZN(n58));
   AOI22_X1 U307 (.A1(FE_OFN29_n171),
	.A2(RS2[2]),
	.B1(FE_OFN92_n170),
	.B2(IR_IN[22]),
	.ZN(n193));
   INV_X1 U308 (.A(n176),
	.ZN(n90));
   AOI22_X1 U309 (.A1(IR_IN[5]),
	.A2(FE_OFN92_n170),
	.B1(OPCODE[5]),
	.B2(FE_OFN29_n171),
	.ZN(n176));
   INV_X1 U310 (.A(n186),
	.ZN(n72));
   AOI22_X1 U311 (.A1(FE_OFN29_n171),
	.A2(RS1[0]),
	.B1(FE_OFN92_n170),
	.B2(IR_IN[15]),
	.ZN(n186));
   INV_X1 U312 (.A(n191),
	.ZN(n62));
   AOI22_X1 U313 (.A1(FE_OFN29_n171),
	.A2(RS2[0]),
	.B1(FE_OFN92_n170),
	.B2(IR_IN[20]),
	.ZN(n191));
   INV_X1 U314 (.A(n187),
	.ZN(n70));
   AOI22_X1 U315 (.A1(FE_OFN29_n171),
	.A2(RS1[1]),
	.B1(FE_OFN92_n170),
	.B2(IR_IN[16]),
	.ZN(n187));
   INV_X1 U316 (.A(n192),
	.ZN(n60));
   AOI22_X1 U317 (.A1(FE_OFN29_n171),
	.A2(RS2[1]),
	.B1(FE_OFN92_n170),
	.B2(IR_IN[21]),
	.ZN(n192));
   INV_X1 U318 (.A(n190),
	.ZN(n64));
   AOI22_X1 U319 (.A1(FE_OFN29_n171),
	.A2(RS1[4]),
	.B1(FE_OFN92_n170),
	.B2(IR_IN[19]),
	.ZN(n190));
   INV_X1 U320 (.A(n195),
	.ZN(n54));
   AOI22_X1 U321 (.A1(FE_OFN29_n171),
	.A2(RS2[4]),
	.B1(FE_OFN92_n170),
	.B2(IR_IN[24]),
	.ZN(n195));
   INV_X1 U322 (.A(n189),
	.ZN(n66));
   AOI22_X1 U323 (.A1(FE_OFN29_n171),
	.A2(RS1[3]),
	.B1(FE_OFN92_n170),
	.B2(IR_IN[18]),
	.ZN(n189));
   INV_X1 U324 (.A(n194),
	.ZN(n56));
   AOI22_X1 U325 (.A1(FE_OFN29_n171),
	.A2(RS2[3]),
	.B1(FE_OFN92_n170),
	.B2(IR_IN[23]),
	.ZN(n194));
   INV_X1 U326 (.A(n175),
	.ZN(n91));
   AOI22_X1 U327 (.A1(IR_IN[4]),
	.A2(FE_OFN92_n170),
	.B1(OPCODE[4]),
	.B2(FE_OFN29_n171),
	.ZN(n175));
   INV_X1 U328 (.A(n174),
	.ZN(n92));
   AOI22_X1 U329 (.A1(IR_IN[3]),
	.A2(FE_OFN92_n170),
	.B1(OPCODE[3]),
	.B2(FE_OFN29_n171),
	.ZN(n174));
   INV_X1 U330 (.A(n178),
	.ZN(n88));
   AOI22_X1 U331 (.A1(FE_OFN29_n171),
	.A2(RD[0]),
	.B1(FE_OFN92_n170),
	.B2(IR_IN[7]),
	.ZN(n178));
   INV_X1 U332 (.A(n179),
	.ZN(n86));
   AOI22_X1 U333 (.A1(FE_OFN29_n171),
	.A2(RD[1]),
	.B1(FE_OFN92_n170),
	.B2(IR_IN[8]),
	.ZN(n179));
   INV_X1 U334 (.A(n180),
	.ZN(n84));
   AOI22_X1 U335 (.A1(FE_OFN29_n171),
	.A2(RD[2]),
	.B1(FE_OFN92_n170),
	.B2(IR_IN[9]),
	.ZN(n180));
   INV_X1 U336 (.A(n181),
	.ZN(n82));
   AOI22_X1 U337 (.A1(FE_OFN29_n171),
	.A2(RD[3]),
	.B1(FE_OFN92_n170),
	.B2(IR_IN[10]),
	.ZN(n181));
   INV_X1 U338 (.A(n182),
	.ZN(n80));
   AOI22_X1 U339 (.A1(FE_OFN29_n171),
	.A2(RD[4]),
	.B1(FE_OFN92_n170),
	.B2(IR_IN[11]),
	.ZN(n182));
   INV_X1 U340 (.A(n183),
	.ZN(n78));
   AOI22_X1 U341 (.A1(FE_OFN29_n171),
	.A2(FUNC3[0]),
	.B1(FE_OFN92_n170),
	.B2(IR_IN[12]),
	.ZN(n183));
   INV_X1 U342 (.A(n177),
	.ZN(n89));
   AOI22_X1 U343 (.A1(IR_IN[6]),
	.A2(FE_OFN92_n170),
	.B1(OPCODE[6]),
	.B2(FE_OFN29_n171),
	.ZN(n177));
   INV_X1 U344 (.A(n202),
	.ZN(n40));
   AOI22_X1 U345 (.A1(FE_OFN29_n171),
	.A2(IMM[31]),
	.B1(FE_OFN92_n170),
	.B2(IR_IN[31]),
	.ZN(n202));
   NOR2_X1 U346 (.A1(FE_OFN35_n205),
	.A2(rst),
	.ZN(n204));
   NOR2_X1 U347 (.A1(rst),
	.A2(en),
	.ZN(n205));
   INV_X1 U348 (.A(EXE_MEM_IN[20]),
	.ZN(n362));
   INV_X1 U349 (.A(EXE_MEM_IN[28]),
	.ZN(n165));
   INV_X1 U350 (.A(EXE_MEM_IN[24]),
	.ZN(n250));
   INV_X1 U351 (.A(EXE_MEM_IN[17]),
	.ZN(n365));
   INV_X1 U352 (.A(EXE_MEM_IN[16]),
	.ZN(n366));
   INV_X1 U353 (.A(EXE_MEM_IN[13]),
	.ZN(n369));
   INV_X1 U354 (.A(EXE_MEM_IN[12]),
	.ZN(n370));
   INV_X1 U355 (.A(EXE_MEM_IN[9]),
	.ZN(n373));
   INV_X1 U356 (.A(EXE_MEM_IN[8]),
	.ZN(n374));
   INV_X1 U357 (.A(EXE_MEM_IN[5]),
	.ZN(n377));
   INV_X1 U358 (.A(EXE_MEM_IN[4]),
	.ZN(n378));
   INV_X1 U359 (.A(EXE_MEM_IN[1]),
	.ZN(n381));
   INV_X1 U360 (.A(EXE_MEM_IN[0]),
	.ZN(n382));
   INV_X1 U361 (.A(n207),
	.ZN(n159));
   AOI22_X1 U362 (.A1(PC_IN[2]),
	.A2(FE_OFN93_n204),
	.B1(PC_OUT[2]),
	.B2(FE_OFN35_n205),
	.ZN(n207));
   INV_X1 U363 (.A(n203),
	.ZN(n161));
   AOI22_X1 U364 (.A1(PC_IN[0]),
	.A2(FE_OFN93_n204),
	.B1(PC_OUT[0]),
	.B2(FE_OFN35_n205),
	.ZN(n203));
   INV_X1 U365 (.A(n208),
	.ZN(n158));
   AOI22_X1 U366 (.A1(PC_IN[3]),
	.A2(FE_OFN93_n204),
	.B1(PC_OUT[3]),
	.B2(FE_OFN35_n205),
	.ZN(n208));
   INV_X1 U367 (.A(n209),
	.ZN(n157));
   AOI22_X1 U368 (.A1(PC_IN[4]),
	.A2(FE_OFN93_n204),
	.B1(PC_OUT[4]),
	.B2(FE_OFN35_n205),
	.ZN(n209));
   INV_X1 U369 (.A(n210),
	.ZN(n156));
   AOI22_X1 U370 (.A1(PC_IN[5]),
	.A2(FE_OFN93_n204),
	.B1(PC_OUT[5]),
	.B2(FE_OFN35_n205),
	.ZN(n210));
   INV_X1 U371 (.A(n211),
	.ZN(n155));
   AOI22_X1 U372 (.A1(PC_IN[6]),
	.A2(FE_OFN93_n204),
	.B1(PC_OUT[6]),
	.B2(FE_OFN35_n205),
	.ZN(n211));
   INV_X1 U373 (.A(n212),
	.ZN(n154));
   AOI22_X1 U374 (.A1(PC_IN[7]),
	.A2(FE_OFN93_n204),
	.B1(PC_OUT[7]),
	.B2(FE_OFN35_n205),
	.ZN(n212));
   INV_X1 U375 (.A(n213),
	.ZN(n153));
   AOI22_X1 U376 (.A1(PC_IN[8]),
	.A2(FE_OFN93_n204),
	.B1(PC_OUT[8]),
	.B2(FE_OFN35_n205),
	.ZN(n213));
   INV_X1 U377 (.A(n214),
	.ZN(n152));
   AOI22_X1 U378 (.A1(PC_IN[9]),
	.A2(FE_OFN93_n204),
	.B1(PC_OUT[9]),
	.B2(FE_OFN35_n205),
	.ZN(n214));
   INV_X1 U379 (.A(n215),
	.ZN(n151));
   AOI22_X1 U380 (.A1(PC_IN[10]),
	.A2(FE_OFN93_n204),
	.B1(PC_OUT[10]),
	.B2(FE_OFN35_n205),
	.ZN(n215));
   INV_X1 U381 (.A(n216),
	.ZN(n150));
   AOI22_X1 U382 (.A1(PC_IN[11]),
	.A2(FE_OFN93_n204),
	.B1(PC_OUT[11]),
	.B2(FE_OFN35_n205),
	.ZN(n216));
   INV_X1 U383 (.A(n217),
	.ZN(n149));
   AOI22_X1 U384 (.A1(PC_IN[12]),
	.A2(FE_OFN93_n204),
	.B1(PC_OUT[12]),
	.B2(FE_OFN35_n205),
	.ZN(n217));
   INV_X1 U385 (.A(n218),
	.ZN(n148));
   AOI22_X1 U386 (.A1(PC_IN[13]),
	.A2(FE_OFN93_n204),
	.B1(PC_OUT[13]),
	.B2(FE_OFN35_n205),
	.ZN(n218));
   INV_X1 U387 (.A(n219),
	.ZN(n147));
   AOI22_X1 U388 (.A1(PC_IN[14]),
	.A2(FE_OFN93_n204),
	.B1(PC_OUT[14]),
	.B2(FE_OFN35_n205),
	.ZN(n219));
   INV_X1 U389 (.A(n220),
	.ZN(n146));
   AOI22_X1 U390 (.A1(PC_IN[15]),
	.A2(FE_OFN93_n204),
	.B1(PC_OUT[15]),
	.B2(FE_OFN35_n205),
	.ZN(n220));
   INV_X1 U391 (.A(n221),
	.ZN(n145));
   AOI22_X1 U392 (.A1(PC_IN[16]),
	.A2(FE_OFN93_n204),
	.B1(PC_OUT[16]),
	.B2(FE_OFN35_n205),
	.ZN(n221));
   INV_X1 U393 (.A(n222),
	.ZN(n144));
   AOI22_X1 U394 (.A1(PC_IN[17]),
	.A2(FE_OFN93_n204),
	.B1(PC_OUT[17]),
	.B2(FE_OFN35_n205),
	.ZN(n222));
   INV_X1 U427 (.A(n223),
	.ZN(n143));
   AOI22_X1 U429 (.A1(PC_IN[18]),
	.A2(FE_OFN93_n204),
	.B1(PC_OUT[18]),
	.B2(FE_OFN35_n205),
	.ZN(n223));
   INV_X1 U430 (.A(n224),
	.ZN(n142));
   AOI22_X1 U431 (.A1(PC_IN[19]),
	.A2(FE_OFN93_n204),
	.B1(PC_OUT[19]),
	.B2(FE_OFN35_n205),
	.ZN(n224));
   INV_X1 U432 (.A(n225),
	.ZN(n141));
   AOI22_X1 U433 (.A1(PC_IN[20]),
	.A2(FE_OFN93_n204),
	.B1(PC_OUT[20]),
	.B2(FE_OFN35_n205),
	.ZN(n225));
   INV_X1 U434 (.A(n226),
	.ZN(n140));
   AOI22_X1 U435 (.A1(PC_IN[21]),
	.A2(FE_OFN93_n204),
	.B1(PC_OUT[21]),
	.B2(FE_OFN35_n205),
	.ZN(n226));
   INV_X1 U436 (.A(n227),
	.ZN(n139));
   AOI22_X1 U437 (.A1(PC_IN[22]),
	.A2(FE_OFN93_n204),
	.B1(PC_OUT[22]),
	.B2(FE_OFN35_n205),
	.ZN(n227));
   INV_X1 U438 (.A(n228),
	.ZN(n138));
   AOI22_X1 U439 (.A1(PC_IN[23]),
	.A2(FE_OFN93_n204),
	.B1(PC_OUT[23]),
	.B2(FE_OFN35_n205),
	.ZN(n228));
   INV_X1 U440 (.A(n229),
	.ZN(n137));
   AOI22_X1 U441 (.A1(PC_IN[24]),
	.A2(FE_OFN93_n204),
	.B1(PC_OUT[24]),
	.B2(FE_OFN35_n205),
	.ZN(n229));
   INV_X1 U442 (.A(n230),
	.ZN(n136));
   AOI22_X1 U443 (.A1(PC_IN[25]),
	.A2(FE_OFN93_n204),
	.B1(PC_OUT[25]),
	.B2(FE_OFN35_n205),
	.ZN(n230));
   INV_X1 U444 (.A(n231),
	.ZN(n135));
   AOI22_X1 U445 (.A1(PC_IN[26]),
	.A2(FE_OFN93_n204),
	.B1(PC_OUT[26]),
	.B2(FE_OFN35_n205),
	.ZN(n231));
   INV_X1 U446 (.A(n232),
	.ZN(n134));
   AOI22_X1 U447 (.A1(PC_IN[27]),
	.A2(FE_OFN93_n204),
	.B1(PC_OUT[27]),
	.B2(FE_OFN35_n205),
	.ZN(n232));
   INV_X1 U448 (.A(n233),
	.ZN(n133));
   AOI22_X1 U449 (.A1(PC_IN[28]),
	.A2(FE_OFN93_n204),
	.B1(PC_OUT[28]),
	.B2(FE_OFN35_n205),
	.ZN(n233));
   INV_X1 U450 (.A(n234),
	.ZN(n132));
   AOI22_X1 U451 (.A1(PC_IN[29]),
	.A2(FE_OFN93_n204),
	.B1(PC_OUT[29]),
	.B2(FE_OFN35_n205),
	.ZN(n234));
   INV_X1 U452 (.A(n235),
	.ZN(n131));
   AOI22_X1 U453 (.A1(PC_IN[30]),
	.A2(FE_OFN93_n204),
	.B1(PC_OUT[30]),
	.B2(FE_OFN35_n205),
	.ZN(n235));
   INV_X1 U454 (.A(n236),
	.ZN(n130));
   AOI22_X1 U455 (.A1(PC_IN[31]),
	.A2(FE_OFN93_n204),
	.B1(PC_OUT[31]),
	.B2(FE_OFN35_n205),
	.ZN(n236));
   INV_X1 U456 (.A(n206),
	.ZN(n160));
   AOI22_X1 U457 (.A1(PC_IN[1]),
	.A2(FE_OFN93_n204),
	.B1(PC_OUT[1]),
	.B2(FE_OFN35_n205),
	.ZN(n206));
   AOI22_X1 U458 (.A1(IR_IN[0]),
	.A2(FE_OFN92_n170),
	.B1(n7),
	.B2(FE_OFN29_n171),
	.ZN(n169));
endmodule

module alu_N32_DW01_add_0 (
	A, 
	B, 
	CI, 
	SUM, 
	CO);
   input [31:0] A;
   input [31:0] B;
   input CI;
   output [31:0] SUM;
   output CO;

   // Internal wires
   wire n3;
   wire n4;
   wire n5;
   wire n6;
   wire n8;
   wire n11;
   wire n12;
   wire n27;
   wire n33;
   wire n35;
   wire n36;
   wire n39;
   wire n43;
   wire n49;
   wire n51;
   wire n52;
   wire n54;
   wire n55;
   wire n56;
   wire n57;
   wire n58;
   wire n59;
   wire n60;
   wire n63;
   wire n64;
   wire n65;
   wire n66;
   wire n67;
   wire n68;
   wire n69;
   wire n70;
   wire n71;
   wire n72;
   wire n73;
   wire n74;
   wire n75;
   wire n76;
   wire n77;
   wire n78;
   wire n79;
   wire n80;
   wire n81;
   wire n82;
   wire n83;
   wire n84;
   wire n85;
   wire n86;
   wire n87;
   wire n88;
   wire n89;
   wire n90;
   wire n91;
   wire n92;
   wire n93;
   wire n94;
   wire n95;
   wire n96;
   wire n97;
   wire n100;
   wire n102;
   wire n103;
   wire n105;
   wire n106;
   wire n107;
   wire n108;
   wire n109;
   wire n110;
   wire n111;
   wire n112;
   wire n114;
   wire n115;
   wire n116;
   wire n117;
   wire n119;
   wire n121;
   wire n122;
   wire n123;
   wire n124;
   wire n125;
   wire n126;
   wire n127;
   wire n128;
   wire n129;
   wire n130;
   wire n131;
   wire n133;
   wire n134;
   wire n135;
   wire n136;
   wire n137;
   wire n140;
   wire n141;
   wire n142;
   wire n143;
   wire n144;
   wire n145;
   wire n146;
   wire n147;
   wire n148;
   wire n149;
   wire n150;
   wire n151;
   wire n152;
   wire n153;
   wire n154;
   wire n155;
   wire n156;
   wire n157;
   wire n158;
   wire n159;
   wire n160;
   wire n161;
   wire n162;
   wire n163;
   wire n164;
   wire n167;
   wire n168;
   wire n169;
   wire n170;
   wire n171;
   wire n172;
   wire n173;
   wire n174;
   wire n175;
   wire n176;
   wire n177;
   wire n178;
   wire n179;
   wire n180;
   wire n181;
   wire n182;
   wire n183;
   wire n184;
   wire n185;
   wire n186;
   wire n187;
   wire n188;
   wire n189;
   wire n190;
   wire n191;
   wire n192;
   wire n194;
   wire n195;
   wire n196;
   wire n197;
   wire n198;
   wire n199;
   wire n200;
   wire n201;
   wire n202;
   wire n203;
   wire n204;
   wire n205;
   wire n206;
   wire n207;
   wire [30:2] carry;

   NAND3_X1 U3 (.A1(n92),
	.A2(n91),
	.A3(n93),
	.ZN(n3));
   NAND2_X1 U4 (.A1(carry[3]),
	.A2(A[3]),
	.ZN(n4));
   NAND2_X1 U5 (.A1(n55),
	.A2(B[8]),
	.ZN(n5));
   NAND2_X1 U6 (.A1(n57),
	.A2(A[15]),
	.ZN(n6));
   NAND3_X1 U8 (.A1(n6),
	.A2(n80),
	.A3(n81),
	.ZN(n8));
   NAND2_X1 U11 (.A1(carry[21]),
	.A2(A[21]),
	.ZN(n11));
   NAND2_X1 U12 (.A1(n164),
	.A2(B[3]),
	.ZN(n12));
   NAND3_X1 U27 (.A1(n69),
	.A2(n68),
	.A3(n70),
	.ZN(n27));
   NAND2_X1 U33 (.A1(n164),
	.A2(B[3]),
	.ZN(n33));
   NAND3_X1 U35 (.A1(n12),
	.A2(n4),
	.A3(n194),
	.ZN(n35));
   NAND3_X1 U36 (.A1(n169),
	.A2(n168),
	.A3(n170),
	.ZN(n36));
   NAND2_X1 U39 (.A1(n59),
	.A2(B[1]),
	.ZN(n39));
   NAND2_X1 U43 (.A1(n59),
	.A2(B[1]),
	.ZN(n43));
   XOR2_X1 U47 (.A(B[31]),
	.B(A[31]),
	.Z(n129));
   NAND3_X1 U50 (.A1(n122),
	.A2(n123),
	.A3(n124),
	.ZN(n49));
   NAND3_X1 U52 (.A1(n95),
	.A2(n97),
	.A3(n96),
	.ZN(n51));
   NAND3_X1 U53 (.A1(n88),
	.A2(n87),
	.A3(n89),
	.ZN(n52));
   NAND3_X1 U55 (.A1(n154),
	.A2(n153),
	.A3(n155),
	.ZN(n54));
   NAND3_X1 U56 (.A1(n162),
	.A2(n161),
	.A3(n163),
	.ZN(n55));
   NAND3_X1 U57 (.A1(n5),
	.A2(n131),
	.A3(n133),
	.ZN(n56));
   NAND3_X1 U58 (.A1(n176),
	.A2(n178),
	.A3(n177),
	.ZN(n57));
   NAND3_X1 U59 (.A1(n11),
	.A2(n150),
	.A3(n151),
	.ZN(n58));
   AND2_X1 U60 (.A1(B[0]),
	.A2(A[0]),
	.ZN(n59));
   NAND3_X1 U61 (.A1(n197),
	.A2(n196),
	.A3(n198),
	.ZN(n60));
   NAND3_X1 U64 (.A1(n204),
	.A2(n205),
	.A3(n206),
	.ZN(n63));
   NAND3_X1 U65 (.A1(n127),
	.A2(n126),
	.A3(n128),
	.ZN(n64));
   NAND3_X1 U66 (.A1(n201),
	.A2(n200),
	.A3(n202),
	.ZN(n65));
   NAND3_X1 U67 (.A1(n110),
	.A2(n111),
	.A3(n112),
	.ZN(n66));
   XOR2_X1 U68 (.A(A[16]),
	.B(B[16]),
	.Z(n67));
   XOR2_X1 U69 (.A(n8),
	.B(n67),
	.Z(SUM[16]));
   NAND2_X1 U70 (.A1(carry[16]),
	.A2(A[16]),
	.ZN(n68));
   NAND2_X1 U71 (.A1(n8),
	.A2(B[16]),
	.ZN(n69));
   NAND2_X1 U72 (.A1(A[16]),
	.A2(B[16]),
	.ZN(n70));
   NAND3_X1 U73 (.A1(n69),
	.A2(n70),
	.A3(n68),
	.ZN(carry[17]));
   NAND3_X1 U74 (.A1(n173),
	.A2(n174),
	.A3(n172),
	.ZN(n71));
   XOR2_X1 U75 (.A(A[25]),
	.B(B[25]),
	.Z(n72));
   XOR2_X1 U76 (.A(n71),
	.B(n72),
	.Z(SUM[25]));
   NAND2_X1 U77 (.A1(n71),
	.A2(A[25]),
	.ZN(n73));
   NAND2_X1 U78 (.A1(carry[25]),
	.A2(B[25]),
	.ZN(n74));
   NAND2_X1 U79 (.A1(A[25]),
	.A2(B[25]),
	.ZN(n75));
   NAND3_X1 U80 (.A1(n73),
	.A2(n74),
	.A3(n75),
	.ZN(carry[26]));
   NAND3_X1 U81 (.A1(n91),
	.A2(n92),
	.A3(n93),
	.ZN(n76));
   AND3_X1 U82 (.A1(n116),
	.A2(n115),
	.A3(n117),
	.ZN(n77));
   XNOR2_X1 U83 (.A(n77),
	.B(n129),
	.ZN(SUM[31]));
   XOR2_X1 U84 (.A(A[15]),
	.B(B[15]),
	.Z(n78));
   XOR2_X1 U85 (.A(n57),
	.B(n78),
	.Z(SUM[15]));
   NAND2_X1 U86 (.A1(n57),
	.A2(A[15]),
	.ZN(n79));
   NAND2_X1 U87 (.A1(carry[15]),
	.A2(B[15]),
	.ZN(n80));
   NAND2_X1 U88 (.A1(A[15]),
	.A2(B[15]),
	.ZN(n81));
   NAND3_X1 U89 (.A1(n79),
	.A2(n80),
	.A3(n81),
	.ZN(carry[16]));
   XOR2_X1 U90 (.A(A[13]),
	.B(B[13]),
	.Z(n82));
   XOR2_X1 U91 (.A(n65),
	.B(n82),
	.Z(SUM[13]));
   NAND2_X1 U92 (.A1(n65),
	.A2(A[13]),
	.ZN(n83));
   NAND2_X1 U93 (.A1(n65),
	.A2(B[13]),
	.ZN(n84));
   NAND2_X1 U94 (.A1(A[13]),
	.A2(B[13]),
	.ZN(n85));
   NAND3_X1 U95 (.A1(n84),
	.A2(n83),
	.A3(n85),
	.ZN(carry[14]));
   XOR2_X1 U96 (.A(A[19]),
	.B(B[19]),
	.Z(n86));
   XOR2_X1 U97 (.A(carry[19]),
	.B(n86),
	.Z(SUM[19]));
   NAND2_X1 U98 (.A1(n64),
	.A2(A[19]),
	.ZN(n87));
   NAND2_X1 U99 (.A1(carry[19]),
	.A2(B[19]),
	.ZN(n88));
   NAND2_X1 U100 (.A1(A[19]),
	.A2(B[19]),
	.ZN(n89));
   XOR2_X1 U102 (.A(A[29]),
	.B(B[29]),
	.Z(n90));
   XOR2_X1 U103 (.A(n60),
	.B(n90),
	.Z(SUM[29]));
   NAND2_X1 U104 (.A1(n60),
	.A2(A[29]),
	.ZN(n91));
   NAND2_X1 U105 (.A1(n60),
	.A2(B[29]),
	.ZN(n92));
   NAND2_X1 U106 (.A1(A[29]),
	.A2(B[29]),
	.ZN(n93));
   XOR2_X1 U108 (.A(A[11]),
	.B(B[11]),
	.Z(n94));
   XOR2_X1 U109 (.A(n63),
	.B(n94),
	.Z(SUM[11]));
   NAND2_X1 U110 (.A1(n63),
	.A2(A[11]),
	.ZN(n95));
   NAND2_X1 U111 (.A1(n63),
	.A2(B[11]),
	.ZN(n96));
   NAND2_X1 U112 (.A1(A[11]),
	.A2(B[11]),
	.ZN(n97));
   NAND3_X1 U113 (.A1(n96),
	.A2(n95),
	.A3(n97),
	.ZN(carry[12]));
   NAND3_X1 U116 (.A1(n149),
	.A2(n150),
	.A3(n151),
	.ZN(n100));
   NAND3_X1 U118 (.A1(n33),
	.A2(n4),
	.A3(n194),
	.ZN(n102));
   NAND3_X1 U119 (.A1(n136),
	.A2(n135),
	.A3(n137),
	.ZN(n103));
   XOR2_X1 U121 (.A(A[26]),
	.B(B[26]),
	.Z(n105));
   XOR2_X1 U122 (.A(carry[26]),
	.B(n105),
	.Z(SUM[26]));
   NAND2_X1 U123 (.A1(carry[26]),
	.A2(A[26]),
	.ZN(n106));
   NAND2_X1 U124 (.A1(carry[26]),
	.A2(B[26]),
	.ZN(n107));
   NAND2_X1 U125 (.A1(A[26]),
	.A2(B[26]),
	.ZN(n108));
   NAND3_X1 U126 (.A1(n106),
	.A2(n107),
	.A3(n108),
	.ZN(carry[27]));
   XOR2_X1 U127 (.A(A[9]),
	.B(B[9]),
	.Z(n109));
   XOR2_X1 U128 (.A(carry[9]),
	.B(n109),
	.Z(SUM[9]));
   NAND2_X1 U129 (.A1(n56),
	.A2(A[9]),
	.ZN(n110));
   NAND2_X1 U130 (.A1(n56),
	.A2(B[9]),
	.ZN(n111));
   NAND2_X1 U131 (.A1(A[9]),
	.A2(B[9]),
	.ZN(n112));
   XOR2_X1 U134 (.A(A[30]),
	.B(B[30]),
	.Z(n114));
   XOR2_X1 U135 (.A(n76),
	.B(n114),
	.Z(SUM[30]));
   NAND2_X1 U136 (.A1(n3),
	.A2(A[30]),
	.ZN(n115));
   NAND2_X1 U137 (.A1(n3),
	.A2(B[30]),
	.ZN(n116));
   NAND2_X1 U138 (.A1(A[30]),
	.A2(B[30]),
	.ZN(n117));
   NAND2_X1 U140 (.A1(A[2]),
	.A2(B[2]),
	.ZN(n119));
   XOR2_X1 U142 (.A(A[17]),
	.B(B[17]),
	.Z(n121));
   XOR2_X1 U143 (.A(carry[17]),
	.B(n121),
	.Z(SUM[17]));
   NAND2_X1 U144 (.A1(carry[17]),
	.A2(A[17]),
	.ZN(n122));
   NAND2_X1 U145 (.A1(n27),
	.A2(B[17]),
	.ZN(n123));
   NAND2_X1 U146 (.A1(A[17]),
	.A2(B[17]),
	.ZN(n124));
   XOR2_X1 U148 (.A(B[18]),
	.B(A[18]),
	.Z(n125));
   XOR2_X1 U149 (.A(n49),
	.B(n125),
	.Z(SUM[18]));
   NAND2_X1 U150 (.A1(n49),
	.A2(B[18]),
	.ZN(n126));
   NAND2_X1 U151 (.A1(n49),
	.A2(A[18]),
	.ZN(n127));
   NAND2_X1 U152 (.A1(B[18]),
	.A2(A[18]),
	.ZN(n128));
   NAND3_X1 U153 (.A1(n127),
	.A2(n128),
	.A3(n126),
	.ZN(carry[19]));
   XOR2_X1 U154 (.A(A[8]),
	.B(B[8]),
	.Z(n130));
   XOR2_X1 U155 (.A(n55),
	.B(n130),
	.Z(SUM[8]));
   NAND2_X1 U156 (.A1(n55),
	.A2(A[8]),
	.ZN(n131));
   NAND2_X1 U158 (.A1(A[8]),
	.A2(B[8]),
	.ZN(n133));
   NAND3_X1 U159 (.A1(n131),
	.A2(n5),
	.A3(n133),
	.ZN(carry[9]));
   XOR2_X1 U160 (.A(B[4]),
	.B(A[4]),
	.Z(n134));
   XOR2_X1 U161 (.A(n35),
	.B(n134),
	.Z(SUM[4]));
   NAND2_X1 U162 (.A1(n102),
	.A2(B[4]),
	.ZN(n135));
   NAND2_X1 U163 (.A1(n35),
	.A2(A[4]),
	.ZN(n136));
   NAND2_X1 U164 (.A1(B[4]),
	.A2(A[4]),
	.ZN(n137));
   NAND3_X1 U165 (.A1(n136),
	.A2(n137),
	.A3(n135),
	.ZN(carry[5]));
   XOR2_X1 U168 (.A(A[20]),
	.B(B[20]),
	.Z(n140));
   XOR2_X1 U169 (.A(n52),
	.B(n140),
	.Z(SUM[20]));
   NAND2_X1 U170 (.A1(n52),
	.A2(A[20]),
	.ZN(n141));
   NAND2_X1 U171 (.A1(n52),
	.A2(B[20]),
	.ZN(n142));
   NAND2_X1 U172 (.A1(A[20]),
	.A2(B[20]),
	.ZN(n143));
   NAND3_X1 U173 (.A1(n142),
	.A2(n141),
	.A3(n143),
	.ZN(carry[21]));
   XOR2_X1 U174 (.A(A[5]),
	.B(B[5]),
	.Z(n144));
   XOR2_X1 U175 (.A(carry[5]),
	.B(n144),
	.Z(SUM[5]));
   NAND2_X1 U176 (.A1(n103),
	.A2(A[5]),
	.ZN(n145));
   NAND2_X1 U177 (.A1(carry[5]),
	.A2(B[5]),
	.ZN(n146));
   NAND2_X1 U178 (.A1(A[5]),
	.A2(B[5]),
	.ZN(n147));
   NAND3_X1 U179 (.A1(n146),
	.A2(n145),
	.A3(n147),
	.ZN(carry[6]));
   XOR2_X1 U180 (.A(A[21]),
	.B(B[21]),
	.Z(n148));
   XOR2_X1 U181 (.A(carry[21]),
	.B(n148),
	.Z(SUM[21]));
   NAND2_X1 U182 (.A1(carry[21]),
	.A2(A[21]),
	.ZN(n149));
   NAND2_X1 U183 (.A1(carry[21]),
	.A2(B[21]),
	.ZN(n150));
   NAND2_X1 U184 (.A1(A[21]),
	.A2(B[21]),
	.ZN(n151));
   XOR2_X1 U186 (.A(A[6]),
	.B(B[6]),
	.Z(n152));
   XOR2_X1 U187 (.A(carry[6]),
	.B(n152),
	.Z(SUM[6]));
   NAND2_X1 U188 (.A1(carry[6]),
	.A2(A[6]),
	.ZN(n153));
   NAND2_X1 U189 (.A1(carry[6]),
	.A2(B[6]),
	.ZN(n154));
   NAND2_X1 U190 (.A1(A[6]),
	.A2(B[6]),
	.ZN(n155));
   XOR2_X1 U192 (.A(A[22]),
	.B(B[22]),
	.Z(n156));
   XOR2_X1 U193 (.A(n58),
	.B(n156),
	.Z(SUM[22]));
   NAND2_X1 U194 (.A1(n58),
	.A2(A[22]),
	.ZN(n157));
   NAND2_X1 U195 (.A1(n100),
	.A2(B[22]),
	.ZN(n158));
   NAND2_X1 U196 (.A1(A[22]),
	.A2(B[22]),
	.ZN(n159));
   NAND3_X1 U197 (.A1(n157),
	.A2(n158),
	.A3(n159),
	.ZN(carry[23]));
   XOR2_X1 U198 (.A(A[7]),
	.B(B[7]),
	.Z(n160));
   XOR2_X1 U199 (.A(n54),
	.B(n160),
	.Z(SUM[7]));
   NAND2_X1 U200 (.A1(n54),
	.A2(A[7]),
	.ZN(n161));
   NAND2_X1 U201 (.A1(n54),
	.A2(B[7]),
	.ZN(n162));
   NAND2_X1 U202 (.A1(A[7]),
	.A2(B[7]),
	.ZN(n163));
   NAND3_X1 U204 (.A1(n191),
	.A2(n190),
	.A3(n189),
	.ZN(n164));
   XOR2_X1 U207 (.A(A[23]),
	.B(B[23]),
	.Z(n167));
   XOR2_X1 U208 (.A(carry[23]),
	.B(n167),
	.Z(SUM[23]));
   NAND2_X1 U209 (.A1(carry[23]),
	.A2(A[23]),
	.ZN(n168));
   NAND2_X1 U210 (.A1(carry[23]),
	.A2(B[23]),
	.ZN(n169));
   NAND2_X1 U211 (.A1(A[23]),
	.A2(B[23]),
	.ZN(n170));
   XOR2_X1 U212 (.A(A[24]),
	.B(B[24]),
	.Z(n171));
   XOR2_X1 U213 (.A(n36),
	.B(n171),
	.Z(SUM[24]));
   NAND2_X1 U214 (.A1(n36),
	.A2(A[24]),
	.ZN(n172));
   NAND2_X1 U215 (.A1(n36),
	.A2(B[24]),
	.ZN(n173));
   NAND2_X1 U216 (.A1(A[24]),
	.A2(B[24]),
	.ZN(n174));
   NAND3_X1 U217 (.A1(n173),
	.A2(n172),
	.A3(n174),
	.ZN(carry[25]));
   XOR2_X1 U218 (.A(A[14]),
	.B(B[14]),
	.Z(n175));
   XOR2_X1 U219 (.A(carry[14]),
	.B(n175),
	.Z(SUM[14]));
   NAND2_X1 U220 (.A1(carry[14]),
	.A2(A[14]),
	.ZN(n176));
   NAND2_X1 U221 (.A1(carry[14]),
	.A2(B[14]),
	.ZN(n177));
   NAND2_X1 U222 (.A1(A[14]),
	.A2(B[14]),
	.ZN(n178));
   NAND3_X1 U223 (.A1(n176),
	.A2(n177),
	.A3(n178),
	.ZN(carry[15]));
   NAND3_X1 U224 (.A1(n39),
	.A2(n187),
	.A3(n186),
	.ZN(n179));
   NAND3_X1 U225 (.A1(n186),
	.A2(n187),
	.A3(n39),
	.ZN(n180));
   XOR2_X1 U226 (.A(A[27]),
	.B(B[27]),
	.Z(n181));
   XOR2_X1 U227 (.A(carry[27]),
	.B(n181),
	.Z(SUM[27]));
   NAND2_X1 U228 (.A1(carry[27]),
	.A2(A[27]),
	.ZN(n182));
   NAND2_X1 U229 (.A1(carry[27]),
	.A2(B[27]),
	.ZN(n183));
   NAND2_X1 U230 (.A1(A[27]),
	.A2(B[27]),
	.ZN(n184));
   NAND3_X1 U231 (.A1(n183),
	.A2(n182),
	.A3(n184),
	.ZN(carry[28]));
   XOR2_X1 U232 (.A(A[1]),
	.B(B[1]),
	.Z(n185));
   XOR2_X1 U233 (.A(n185),
	.B(n59),
	.Z(SUM[1]));
   NAND2_X1 U234 (.A1(B[1]),
	.A2(A[1]),
	.ZN(n186));
   NAND2_X1 U235 (.A1(n207),
	.A2(A[1]),
	.ZN(n187));
   NAND3_X1 U236 (.A1(n187),
	.A2(n43),
	.A3(n186),
	.ZN(carry[2]));
   XOR2_X1 U237 (.A(A[2]),
	.B(B[2]),
	.Z(n188));
   XOR2_X1 U238 (.A(n188),
	.B(n180),
	.Z(SUM[2]));
   NAND2_X1 U239 (.A1(A[2]),
	.A2(B[2]),
	.ZN(n189));
   NAND2_X1 U240 (.A1(carry[2]),
	.A2(A[2]),
	.ZN(n190));
   NAND2_X1 U241 (.A1(n179),
	.A2(B[2]),
	.ZN(n191));
   NAND3_X1 U242 (.A1(n191),
	.A2(n190),
	.A3(n119),
	.ZN(carry[3]));
   XOR2_X1 U243 (.A(B[3]),
	.B(A[3]),
	.Z(n192));
   XOR2_X1 U244 (.A(n164),
	.B(n192),
	.Z(SUM[3]));
   NAND2_X1 U246 (.A1(B[3]),
	.A2(A[3]),
	.ZN(n194));
   XOR2_X1 U247 (.A(A[28]),
	.B(B[28]),
	.Z(n195));
   XOR2_X1 U248 (.A(carry[28]),
	.B(n195),
	.Z(SUM[28]));
   NAND2_X1 U249 (.A1(carry[28]),
	.A2(A[28]),
	.ZN(n196));
   NAND2_X1 U250 (.A1(carry[28]),
	.A2(B[28]),
	.ZN(n197));
   NAND2_X1 U251 (.A1(A[28]),
	.A2(B[28]),
	.ZN(n198));
   XOR2_X1 U253 (.A(A[12]),
	.B(B[12]),
	.Z(n199));
   XOR2_X1 U254 (.A(n51),
	.B(n199),
	.Z(SUM[12]));
   NAND2_X1 U255 (.A1(carry[12]),
	.A2(A[12]),
	.ZN(n200));
   NAND2_X1 U256 (.A1(n51),
	.A2(B[12]),
	.ZN(n201));
   NAND2_X1 U257 (.A1(A[12]),
	.A2(B[12]),
	.ZN(n202));
   XOR2_X1 U259 (.A(A[10]),
	.B(B[10]),
	.Z(n203));
   XOR2_X1 U260 (.A(n66),
	.B(n203),
	.Z(SUM[10]));
   NAND2_X1 U261 (.A1(n66),
	.A2(A[10]),
	.ZN(n204));
   NAND2_X1 U262 (.A1(n66),
	.A2(B[10]),
	.ZN(n205));
   NAND2_X1 U263 (.A1(A[10]),
	.A2(B[10]),
	.ZN(n206));
   AND2_X1 U265 (.A1(B[0]),
	.A2(A[0]),
	.ZN(n207));
   XOR2_X1 U266 (.A(B[0]),
	.B(A[0]),
	.Z(SUM[0]));
endmodule

module alu_N32_DW_cmp_0 (
	A, 
	B, 
	TC, 
	GE_LT, 
	GE_GT_EQ, 
	GE_LT_GT_LE, 
	EQ_NE, 
	n188, 
	n33);
   input [31:0] A;
   input [31:0] B;
   input TC;
   input GE_LT;
   input GE_GT_EQ;
   output GE_LT_GT_LE;
   output EQ_NE;
   input n188;
   input n33;

   // Internal wires
   wire FE_RN_2_0;
   wire FE_RN_1_0;
   wire FE_RN_0_0;
   wire FE_OFN129_ALU_OPB_16;
   wire n1311;
   wire n1312;
   wire n1314;
   wire n1315;
   wire n1316;
   wire n1317;
   wire n1318;
   wire n1320;
   wire n1322;
   wire n1323;
   wire n1325;
   wire n1331;
   wire n1332;
   wire n1333;
   wire n1336;
   wire n1338;
   wire n1339;
   wire n1340;
   wire n1341;
   wire n1342;
   wire n1343;
   wire n1344;
   wire n1345;
   wire n1346;
   wire n1347;
   wire n1348;
   wire n1349;
   wire n1351;
   wire n1352;
   wire n1353;
   wire n1354;
   wire n1355;
   wire n1356;
   wire n1357;
   wire n1358;
   wire n1359;
   wire n1360;
   wire n1361;
   wire n1362;
   wire n1363;
   wire n1364;
   wire n1365;
   wire n1366;
   wire n1367;
   wire n1368;
   wire n1369;
   wire n1370;
   wire n1371;
   wire n1372;
   wire n1373;
   wire n1374;
   wire n1375;
   wire n1376;
   wire n1377;
   wire n1378;
   wire n1379;
   wire n1380;
   wire n1381;
   wire n1382;
   wire n1383;
   wire n1384;
   wire n1385;
   wire n1386;
   wire n1387;
   wire n1388;
   wire n1389;
   wire n1390;
   wire n1391;
   wire n1392;
   wire n1393;
   wire n1394;
   wire n1395;
   wire n1396;
   wire n1397;
   wire n1398;
   wire n1399;
   wire n1400;
   wire n1401;
   wire n1402;
   wire n1403;
   wire n1404;
   wire n1405;
   wire n1406;
   wire n1407;
   wire n1408;
   wire n1409;
   wire n1410;
   wire n1411;
   wire n1412;
   wire n1413;
   wire n1414;
   wire n1415;
   wire n1416;
   wire n1417;
   wire n1418;
   wire n1419;
   wire n1420;
   wire n1421;
   wire n1422;
   wire n1423;
   wire n1424;
   wire n1425;
   wire n1426;
   wire n1427;
   wire n1428;
   wire n1429;
   wire n1430;
   wire n1431;
   wire n1432;

   INV_X1 FE_RC_10_0 (.A(n1390),
	.ZN(FE_RN_2_0));
   AOI21_X1 FE_RC_9_0 (.A(n1384),
	.B1(FE_RN_2_0),
	.B2(n1385),
	.ZN(n1376));
   AOI21_X1 FE_RC_8_0 (.A(n1369),
	.B1(n1320),
	.B2(n1370),
	.ZN(n1361));
   AOI21_X1 FE_RC_7_0 (.A(n1357),
	.B1(n1358),
	.B2(n1359),
	.ZN(n1356));
   AOI21_X1 FE_RC_6_0 (.A(n1418),
	.B1(n1316),
	.B2(n1419),
	.ZN(n1417));
   AOI21_X1 FE_RC_5_0 (.A(n1378),
	.B1(n1333),
	.B2(n1379),
	.ZN(n1377));
   AOI21_X1 FE_RC_4_0 (.A(n1363),
	.B1(n1325),
	.B2(n1364),
	.ZN(n1362));
   INV_X1 FE_RC_3_0 (.A(n1406),
	.ZN(FE_RN_1_0));
   AOI21_X1 FE_RC_2_0 (.A(n1400),
	.B1(FE_RN_1_0),
	.B2(n1401),
	.ZN(n1399));
   INV_X1 FE_RC_1_0 (.A(n1430),
	.ZN(FE_RN_0_0));
   AOI21_X1 FE_RC_0_0 (.A(n1424),
	.B1(FE_RN_0_0),
	.B2(n1425),
	.ZN(n1416));
   BUF_X1 FE_OFC129_ALU_OPB_16 (.A(B[16]),
	.Z(FE_OFN129_ALU_OPB_16));
   INV_X1 U655 (.A(n1398),
	.ZN(n1318));
   INV_X1 U657 (.A(n1360),
	.ZN(n1323));
   INV_X1 U659 (.A(n1410),
	.ZN(n1331));
   INV_X1 U660 (.A(n1411),
	.ZN(n1312));
   INV_X1 U661 (.A(A[1]),
	.ZN(n1322));
   INV_X1 U666 (.A(A[10]),
	.ZN(n1314));
   INV_X1 U667 (.A(A[12]),
	.ZN(n1315));
   INV_X1 U668 (.A(A[14]),
	.ZN(n1317));
   INV_X1 U676 (.A(B[25]),
	.ZN(n1347));
   INV_X1 U677 (.A(B[19]),
	.ZN(n1344));
   INV_X1 U678 (.A(B[23]),
	.ZN(n1346));
   INV_X1 U679 (.A(B[9]),
	.ZN(n1353));
   INV_X1 U680 (.A(B[21]),
	.ZN(n1345));
   INV_X1 U681 (.A(A[2]),
	.ZN(n1332));
   INV_X1 U682 (.A(A[8]),
	.ZN(n1339));
   INV_X1 U683 (.A(A[6]),
	.ZN(n1338));
   INV_X1 U684 (.A(A[4]),
	.ZN(n1336));
   INV_X1 U685 (.A(B[5]),
	.ZN(n1351));
   INV_X1 U686 (.A(B[29]),
	.ZN(n1349));
   INV_X1 U687 (.A(B[27]),
	.ZN(n1348));
   INV_X1 U688 (.A(B[7]),
	.ZN(n1352));
   INV_X1 U689 (.A(B[17]),
	.ZN(n1343));
   INV_X1 U690 (.A(n1392),
	.ZN(n1325));
   INV_X1 U691 (.A(n1391),
	.ZN(n1320));
   INV_X1 U692 (.A(n1407),
	.ZN(n1311));
   INV_X1 U693 (.A(n1394),
	.ZN(n1333));
   INV_X1 U694 (.A(n1432),
	.ZN(n1316));
   INV_X1 U695 (.A(B[13]),
	.ZN(n1341));
   INV_X1 U696 (.A(B[11]),
	.ZN(n1340));
   INV_X1 U697 (.A(B[15]),
	.ZN(n1342));
   OAI21_X1 U699 (.A(n1356),
	.B1(n1354),
	.B2(n1355),
	.ZN(GE_LT_GT_LE));
   OAI21_X1 U701 (.A(n1362),
	.B1(n1360),
	.B2(n1361),
	.ZN(n1358));
   OAI21_X1 U703 (.A(n1365),
	.B1(A[21]),
	.B2(n1345),
	.ZN(n1364));
   NAND3_X1 U704 (.A1(n1366),
	.A2(A[20]),
	.A3(B[20]),
	.ZN(n1365));
   OAI21_X1 U705 (.A(n1367),
	.B1(A[23]),
	.B2(n1346),
	.ZN(n1363));
   NAND3_X1 U706 (.A1(n1368),
	.A2(A[22]),
	.A3(B[22]),
	.ZN(n1367));
   OAI21_X1 U708 (.A(n1371),
	.B1(A[17]),
	.B2(n1343),
	.ZN(n1370));
   NAND3_X1 U709 (.A1(n1372),
	.A2(A[16]),
	.A3(FE_OFN129_ALU_OPB_16),
	.ZN(n1371));
   OAI21_X1 U710 (.A(n1373),
	.B1(A[19]),
	.B2(n1344),
	.ZN(n1369));
   NAND3_X1 U711 (.A1(n1374),
	.A2(A[18]),
	.A3(B[18]),
	.ZN(n1373));
   OAI21_X1 U712 (.A(n1377),
	.B1(n1375),
	.B2(n1376),
	.ZN(n1357));
   OAI21_X1 U714 (.A(n1380),
	.B1(A[29]),
	.B2(n1349),
	.ZN(n1379));
   NAND3_X1 U715 (.A1(n1381),
	.A2(A[28]),
	.A3(B[28]),
	.ZN(n1380));
   OAI21_X1 U716 (.A(n1382),
	.B1(B[31]),
	.B2(A[31]),
	.ZN(n1378));
   NAND3_X1 U717 (.A1(n1383),
	.A2(A[30]),
	.A3(B[30]),
	.ZN(n1382));
   OAI21_X1 U719 (.A(n1386),
	.B1(A[25]),
	.B2(n1347),
	.ZN(n1385));
   NAND3_X1 U720 (.A1(n1387),
	.A2(A[24]),
	.A3(B[24]),
	.ZN(n1386));
   OAI21_X1 U721 (.A(n1388),
	.B1(A[27]),
	.B2(n1348),
	.ZN(n1384));
   NAND3_X1 U722 (.A1(n1389),
	.A2(A[26]),
	.A3(B[26]),
	.ZN(n1388));
   NAND3_X1 U723 (.A1(n1359),
	.A2(n1323),
	.A3(n1320),
	.ZN(n1355));
   OAI21_X1 U724 (.A(n1374),
	.B1(B[18]),
	.B2(A[18]),
	.ZN(n1391));
   NAND2_X1 U725 (.A1(A[19]),
	.A2(n1344),
	.ZN(n1374));
   OAI211_X1 U726 (.A(n1366),
	.B(n1325),
	.C1(B[20]),
	.C2(A[20]),
	.ZN(n1360));
   OAI21_X1 U727 (.A(n1368),
	.B1(B[22]),
	.B2(A[22]),
	.ZN(n1392));
   NAND2_X1 U728 (.A1(A[23]),
	.A2(n1346),
	.ZN(n1368));
   NAND2_X1 U729 (.A1(A[21]),
	.A2(n1345),
	.ZN(n1366));
   NOR3_X1 U730 (.A1(n1390),
	.A2(n1375),
	.A3(n1393),
	.ZN(n1359));
   OAI21_X1 U731 (.A(n1387),
	.B1(A[24]),
	.B2(B[24]),
	.ZN(n1393));
   NAND2_X1 U732 (.A1(A[25]),
	.A2(n1347),
	.ZN(n1387));
   OAI211_X1 U733 (.A(n1381),
	.B(n1333),
	.C1(B[28]),
	.C2(A[28]),
	.ZN(n1375));
   OAI21_X1 U734 (.A(n1383),
	.B1(B[30]),
	.B2(A[30]),
	.ZN(n1394));
   NAND2_X1 U735 (.A1(B[31]),
	.A2(A[31]),
	.ZN(n1383));
   NAND2_X1 U736 (.A1(A[29]),
	.A2(n1349),
	.ZN(n1381));
   OAI21_X1 U737 (.A(n1389),
	.B1(B[26]),
	.B2(A[26]),
	.ZN(n1390));
   NAND2_X1 U738 (.A1(A[27]),
	.A2(n1348),
	.ZN(n1389));
   OAI221_X1 U739 (.A(n1318),
	.B1(n1395),
	.B2(n1396),
	.C1(n1396),
	.C2(n1397),
	.ZN(n1354));
   OAI21_X1 U740 (.A(n1372),
	.B1(A[16]),
	.B2(FE_OFN129_ALU_OPB_16),
	.ZN(n1398));
   NAND2_X1 U741 (.A1(A[17]),
	.A2(n1343),
	.ZN(n1372));
   NAND2_X1 U742 (.A1(n1311),
	.A2(n1399),
	.ZN(n1397));
   OAI21_X1 U744 (.A(n1402),
	.B1(A[5]),
	.B2(n1351),
	.ZN(n1401));
   NAND3_X1 U745 (.A1(n1403),
	.A2(n1336),
	.A3(B[4]),
	.ZN(n1402));
   OAI21_X1 U746 (.A(n1404),
	.B1(A[7]),
	.B2(n1352),
	.ZN(n1400));
   NAND3_X1 U747 (.A1(n1405),
	.A2(n1338),
	.A3(B[6]),
	.ZN(n1404));
   AOI211_X1 U748 (.A(n1406),
	.B(n1409),
	.C1(n1408),
	.C2(n1331),
	.ZN(n1407));
   OAI221_X1 U749 (.A(n1403),
	.B1(n1312),
	.B2(n1410),
	.C1(n1336),
	.C2(B[4]),
	.ZN(n1409));
   NAND2_X1 U750 (.A1(A[5]),
	.A2(n1351),
	.ZN(n1403));
   AOI22_X1 U751 (.A1(B[1]),
	.A2(n1322),
	.B1(n1412),
	.B2(B[0]),
	.ZN(n1411));
   AOI21_X1 U752 (.A(A[0]),
	.B1(A[1]),
	.B2(n188),
	.ZN(n1412));
   OAI21_X1 U753 (.A(n1405),
	.B1(B[6]),
	.B2(n1338),
	.ZN(n1406));
   NAND2_X1 U754 (.A1(A[7]),
	.A2(n1352),
	.ZN(n1405));
   OAI21_X1 U755 (.A(n1413),
	.B1(A[3]),
	.B2(B[3]),
	.ZN(n1410));
   NAND3_X1 U756 (.A1(n1414),
	.A2(n1332),
	.A3(n33),
	.ZN(n1413));
   OAI21_X1 U757 (.A(n1414),
	.B1(n1332),
	.B2(n33),
	.ZN(n1408));
   NAND2_X1 U758 (.A1(A[3]),
	.A2(B[3]),
	.ZN(n1414));
   OAI21_X1 U759 (.A(n1417),
	.B1(n1415),
	.B2(n1416),
	.ZN(n1396));
   OAI21_X1 U761 (.A(n1420),
	.B1(A[13]),
	.B2(n1341),
	.ZN(n1419));
   NAND3_X1 U762 (.A1(n1421),
	.A2(n1315),
	.A3(B[12]),
	.ZN(n1420));
   OAI21_X1 U763 (.A(n1422),
	.B1(A[15]),
	.B2(n1342),
	.ZN(n1418));
   NAND3_X1 U764 (.A1(n1423),
	.A2(n1317),
	.A3(B[14]),
	.ZN(n1422));
   OAI21_X1 U766 (.A(n1426),
	.B1(A[9]),
	.B2(n1353),
	.ZN(n1425));
   NAND3_X1 U767 (.A1(n1427),
	.A2(n1339),
	.A3(B[8]),
	.ZN(n1426));
   OAI21_X1 U768 (.A(n1428),
	.B1(A[11]),
	.B2(n1340),
	.ZN(n1424));
   NAND3_X1 U769 (.A1(n1429),
	.A2(n1314),
	.A3(B[10]),
	.ZN(n1428));
   NOR3_X1 U770 (.A1(n1431),
	.A2(n1415),
	.A3(n1430),
	.ZN(n1395));
   OAI21_X1 U771 (.A(n1429),
	.B1(B[10]),
	.B2(n1314),
	.ZN(n1430));
   NAND2_X1 U772 (.A1(A[11]),
	.A2(n1340),
	.ZN(n1429));
   OAI211_X1 U773 (.A(n1421),
	.B(n1316),
	.C1(B[12]),
	.C2(n1315),
	.ZN(n1415));
   OAI21_X1 U774 (.A(n1423),
	.B1(B[14]),
	.B2(n1317),
	.ZN(n1432));
   NAND2_X1 U775 (.A1(A[15]),
	.A2(n1342),
	.ZN(n1423));
   NAND2_X1 U776 (.A1(A[13]),
	.A2(n1341),
	.ZN(n1421));
   OAI21_X1 U777 (.A(n1427),
	.B1(B[8]),
	.B2(n1339),
	.ZN(n1431));
   NAND2_X1 U778 (.A1(A[9]),
	.A2(n1353),
	.ZN(n1427));
endmodule

module alu_N32 (
	OP, 
	ALU_OPA, 
	ALU_OPB, 
	ALU_OUT);
   input [2:0] OP;
   input [31:0] ALU_OPA;
   input [31:0] ALU_OPB;
   output [31:0] ALU_OUT;

   // Internal wires
   wire FE_OFN130_ALU_OPA_0;
   wire FE_OFN128_ALU_OPB_4;
   wire FE_OFN127_ALU_OPA_6;
   wire FE_OFN126_ALU_OPA_8;
   wire FE_OFN125_ALU_OPA_7;
   wire FE_OFN124_ALU_OPA_3;
   wire FE_OFN123_ALU_OPA_5;
   wire FE_OFN122_ALU_OPA_12;
   wire FE_OFN121_ALU_OPA_10;
   wire FE_OFN120_ALU_OPA_14;
   wire FE_OFN119_ALU_OPA_18;
   wire FE_OFN118_ALU_OPA_23;
   wire FE_OFN117_ALU_OPA_24;
   wire FE_OFN116_ALU_OPA_30;
   wire FE_OFN115_ALU_OPB_0;
   wire FE_OFN42_FE_DBTN4_n4;
   wire FE_OFN34_n198;
   wire FE_DBTN15_ALU_OPA_31;
   wire FE_DBTN14_ALU_OPA_30;
   wire FE_DBTN13_ALU_OPA_28;
   wire FE_DBTN12_ALU_OPA_26;
   wire FE_DBTN11_ALU_OPA_24;
   wire FE_DBTN10_ALU_OPA_22;
   wire FE_DBTN9_ALU_OPA_20;
   wire FE_DBTN8_ALU_OPA_18;
   wire FE_DBTN7_ALU_OPA_16;
   wire FE_DBTN6_ALU_OPB_3;
   wire FE_DBTN5_ALU_OPB_0;
   wire FE_DBTN4_n4;
   wire N591;
   wire N613;
   wire N617;
   wire N621;
   wire N625;
   wire N629;
   wire N633;
   wire N637;
   wire N641;
   wire N645;
   wire N649;
   wire N653;
   wire N657;
   wire N661;
   wire N665;
   wire N669;
   wire N671;
   wire N672;
   wire N673;
   wire N674;
   wire N675;
   wire N676;
   wire N677;
   wire N678;
   wire N679;
   wire N680;
   wire N681;
   wire N682;
   wire N683;
   wire N684;
   wire N685;
   wire N686;
   wire N687;
   wire N688;
   wire N689;
   wire N690;
   wire N691;
   wire N692;
   wire N693;
   wire N694;
   wire N695;
   wire N696;
   wire N697;
   wire N698;
   wire N699;
   wire N700;
   wire N701;
   wire N702;
   wire N703;
   wire N335;
   wire N334;
   wire N333;
   wire N332;
   wire N331;
   wire n4;
   wire FE_UNCONNECTED_1;
   wire n9;
   wire n10;
   wire n11;
   wire n12;
   wire n13;
   wire n14;
   wire n15;
   wire n16;
   wire n17;
   wire n18;
   wire n19;
   wire n20;
   wire n21;
   wire n22;
   wire n23;
   wire n24;
   wire n25;
   wire n26;
   wire n27;
   wire n28;
   wire n29;
   wire n30;
   wire n31;
   wire n32;
   wire n33;
   wire n34;
   wire n35;
   wire n36;
   wire n37;
   wire n38;
   wire n39;
   wire n40;
   wire n41;
   wire n42;
   wire n43;
   wire n44;
   wire n45;
   wire n46;
   wire n47;
   wire n48;
   wire n49;
   wire n50;
   wire n51;
   wire n52;
   wire n53;
   wire n54;
   wire n55;
   wire n56;
   wire n57;
   wire n58;
   wire n59;
   wire n60;
   wire n61;
   wire n62;
   wire n63;
   wire n64;
   wire n65;
   wire n66;
   wire n67;
   wire n68;
   wire n69;
   wire n70;
   wire n71;
   wire n72;
   wire n73;
   wire n74;
   wire n75;
   wire n76;
   wire n77;
   wire n78;
   wire n79;
   wire n80;
   wire n81;
   wire n82;
   wire n83;
   wire n84;
   wire n85;
   wire n86;
   wire n87;
   wire n88;
   wire n89;
   wire n90;
   wire n91;
   wire n92;
   wire n93;
   wire n94;
   wire n95;
   wire n96;
   wire n97;
   wire n98;
   wire n99;
   wire n100;
   wire n101;
   wire n102;
   wire n103;
   wire n104;
   wire n105;
   wire n106;
   wire n107;
   wire n108;
   wire n109;
   wire n110;
   wire n111;
   wire n112;
   wire n113;
   wire n114;
   wire n115;
   wire n116;
   wire n117;
   wire n118;
   wire n119;
   wire n120;
   wire n121;
   wire n122;
   wire n123;
   wire n124;
   wire n125;
   wire n126;
   wire n127;
   wire n128;
   wire n129;
   wire n130;
   wire n131;
   wire n133;
   wire n134;
   wire n135;
   wire n137;
   wire n138;
   wire n139;
   wire n140;
   wire n141;
   wire n142;
   wire n143;
   wire n144;
   wire n145;
   wire n146;
   wire n147;
   wire n148;
   wire n149;
   wire n150;
   wire n151;
   wire n152;
   wire n153;
   wire n154;
   wire n170;
   wire n171;
   wire n188;
   wire n189;
   wire n190;
   wire n191;
   wire n192;
   wire n193;
   wire n194;
   wire n198;
   wire n199;
   wire n200;
   wire n201;
   wire n202;
   wire n203;
   wire n204;
   wire n205;
   wire n206;
   wire n207;
   wire n208;
   wire n209;
   wire n210;
   wire n211;
   wire n212;
   wire n213;
   wire n214;
   wire n215;
   wire n216;
   wire n217;
   wire n218;
   wire n219;
   wire n220;
   wire n221;
   wire n222;
   wire n223;
   wire n224;
   wire n225;
   wire n226;
   wire n227;
   wire n228;
   wire n229;
   wire n230;
   wire n231;
   wire n232;
   wire n233;
   wire n234;
   wire n235;
   wire n236;
   wire n237;
   wire n238;
   wire n239;
   wire n240;
   wire n241;
   wire n242;
   wire n243;
   wire n244;
   wire n245;
   wire n246;
   wire n247;
   wire n248;
   wire n249;
   wire n250;
   wire n251;
   wire n252;
   wire n253;
   wire n254;
   wire n255;
   wire n256;
   wire n257;
   wire n258;
   wire n259;
   wire n260;
   wire n261;
   wire n262;
   wire n263;
   wire n264;
   wire n265;
   wire n266;
   wire n267;
   wire n268;
   wire n269;
   wire n270;
   wire n271;
   wire n272;
   wire n273;
   wire n274;
   wire n275;
   wire n276;
   wire n277;
   wire n278;
   wire n279;
   wire n280;
   wire n281;
   wire n282;
   wire n283;
   wire n284;
   wire n285;
   wire n286;
   wire n287;
   wire n288;
   wire n289;
   wire n290;
   wire n291;
   wire n292;
   wire n293;
   wire n294;
   wire n295;
   wire n296;
   wire n297;
   wire n298;
   wire n299;
   wire n300;
   wire n301;
   wire n302;
   wire n303;
   wire n304;
   wire n305;
   wire n307;
   wire n308;
   wire n309;
   wire n310;
   wire n311;
   wire n312;
   wire n313;
   wire n314;
   wire n315;
   wire n316;
   wire n317;
   wire n318;
   wire n319;
   wire n320;
   wire n321;
   wire n322;
   wire n323;
   wire n324;
   wire n325;
   wire n326;
   wire n327;
   wire n328;
   wire n329;
   wire n330;
   wire n331;
   wire n332;
   wire n333;
   wire n334;
   wire n335;
   wire n336;
   wire n337;
   wire n338;
   wire n339;
   wire n340;
   wire n341;
   wire n342;
   wire n343;
   wire n344;
   wire n345;
   wire n346;
   wire n347;
   wire n348;
   wire n349;
   wire n350;
   wire n351;
   wire n352;
   wire n356;
   wire n357;
   wire n358;
   wire n359;
   wire n360;
   wire n361;
   wire n362;
   wire n363;
   wire n364;
   wire n365;
   wire n366;
   wire n367;
   wire n368;
   wire n369;
   wire n370;
   wire n371;
   wire n372;
   wire n373;
   wire n374;
   wire n375;
   wire n376;
   wire n377;
   wire n378;
   wire n379;
   wire n380;
   wire n381;
   wire n382;
   wire n383;
   wire n384;
   wire n386;
   wire n387;
   wire n388;
   wire n389;
   wire n390;
   wire n391;
   wire n392;
   wire n393;
   wire n394;
   wire n395;
   wire n396;
   wire n397;
   wire n398;
   wire n399;
   wire n400;
   wire n401;
   wire n402;
   wire n403;
   wire n404;
   wire n405;
   wire n406;
   wire n407;
   wire n408;
   wire n409;
   wire n410;
   wire n411;
   wire n412;
   wire n413;
   wire n414;
   wire n415;
   wire n417;
   wire n418;
   wire n419;
   wire n420;
   wire n421;
   wire n422;
   wire n423;
   wire n424;
   wire n425;
   wire n426;
   wire n427;
   wire n428;
   wire n429;
   wire n430;
   wire n431;
   wire n432;
   wire n433;
   wire n434;
   wire n435;
   wire n436;
   wire n437;
   wire n438;
   wire n439;
   wire n440;
   wire n441;
   wire n442;
   wire n443;
   wire n444;
   wire n445;
   wire n446;
   wire n447;
   wire n448;
   wire n449;
   wire n450;
   wire n451;
   wire n452;
   wire n453;
   wire n454;
   wire n455;
   wire n456;
   wire n457;
   wire n458;
   wire n459;
   wire n460;
   wire n461;
   wire n462;
   wire n463;
   wire n464;
   wire n465;
   wire n466;
   wire n468;
   wire n469;
   wire n470;
   wire n471;
   wire n472;
   wire n473;
   wire n474;
   wire n475;
   wire n476;
   wire n477;
   wire n478;
   wire n479;
   wire n480;
   wire n481;
   wire n482;
   wire n483;
   wire n484;
   wire n485;
   wire n486;
   wire n487;
   wire n488;
   wire n489;
   wire n490;
   wire n491;
   wire n492;
   wire n493;
   wire n494;
   wire n495;
   wire n496;
   wire n497;
   wire n498;
   wire n499;
   wire n501;
   wire n502;
   wire n503;
   wire n504;
   wire n505;
   wire n506;
   wire n507;
   wire n508;
   wire n509;
   wire n510;
   wire n511;
   wire n512;
   wire n513;
   wire n514;
   wire n515;
   wire n516;
   wire n517;
   wire n518;
   wire n519;
   wire n520;
   wire n521;
   wire n522;
   wire n523;
   wire n524;
   wire n525;
   wire n526;
   wire n527;
   wire n528;
   wire n529;
   wire n530;
   wire n531;
   wire n532;
   wire n533;
   wire n534;
   wire n535;
   wire n536;
   wire n537;
   wire n538;
   wire n539;
   wire n540;
   wire n541;
   wire n542;
   wire n543;
   wire n544;
   wire n545;
   wire n546;
   wire n547;
   wire n548;
   wire n549;
   wire n550;
   wire n551;
   wire n552;
   wire n553;
   wire n554;
   wire n555;
   wire [4:2] r422_carry;

   BUF_X1 FE_OFC130_ALU_OPA_0 (.A(ALU_OPA[0]),
	.Z(FE_OFN130_ALU_OPA_0));
   BUF_X1 FE_OFC128_ALU_OPB_4 (.A(ALU_OPB[4]),
	.Z(FE_OFN128_ALU_OPB_4));
   BUF_X1 FE_OFC127_ALU_OPA_6 (.A(ALU_OPA[6]),
	.Z(FE_OFN127_ALU_OPA_6));
   BUF_X1 FE_OFC126_ALU_OPA_8 (.A(ALU_OPA[8]),
	.Z(FE_OFN126_ALU_OPA_8));
   BUF_X1 FE_OFC125_ALU_OPA_7 (.A(ALU_OPA[7]),
	.Z(FE_OFN125_ALU_OPA_7));
   BUF_X1 FE_OFC124_ALU_OPA_3 (.A(ALU_OPA[3]),
	.Z(FE_OFN124_ALU_OPA_3));
   BUF_X1 FE_OFC123_ALU_OPA_5 (.A(ALU_OPA[5]),
	.Z(FE_OFN123_ALU_OPA_5));
   BUF_X1 FE_OFC122_ALU_OPA_12 (.A(ALU_OPA[12]),
	.Z(FE_OFN122_ALU_OPA_12));
   BUF_X1 FE_OFC121_ALU_OPA_10 (.A(ALU_OPA[10]),
	.Z(FE_OFN121_ALU_OPA_10));
   BUF_X1 FE_OFC120_ALU_OPA_14 (.A(ALU_OPA[14]),
	.Z(FE_OFN120_ALU_OPA_14));
   BUF_X1 FE_OFC119_ALU_OPA_18 (.A(ALU_OPA[18]),
	.Z(FE_OFN119_ALU_OPA_18));
   BUF_X1 FE_OFC118_ALU_OPA_23 (.A(ALU_OPA[23]),
	.Z(FE_OFN118_ALU_OPA_23));
   BUF_X1 FE_OFC117_ALU_OPA_24 (.A(ALU_OPA[24]),
	.Z(FE_OFN117_ALU_OPA_24));
   BUF_X1 FE_OFC116_ALU_OPA_30 (.A(ALU_OPA[30]),
	.Z(FE_OFN116_ALU_OPA_30));
   BUF_X2 FE_OFC115_ALU_OPB_0 (.A(ALU_OPB[0]),
	.Z(FE_OFN115_ALU_OPB_0));
   BUF_X1 FE_OFC42_FE_DBTN4_n4 (.A(FE_DBTN4_n4),
	.Z(FE_OFN42_FE_DBTN4_n4));
   BUF_X2 FE_OFC34_n198 (.A(n198),
	.Z(FE_OFN34_n198));
   INV_X1 FE_DBTC15_ALU_OPA_31 (.A(ALU_OPA[31]),
	.ZN(FE_DBTN15_ALU_OPA_31));
   INV_X1 FE_DBTC14_ALU_OPA_30 (.A(FE_OFN116_ALU_OPA_30),
	.ZN(FE_DBTN14_ALU_OPA_30));
   INV_X1 FE_DBTC13_ALU_OPA_28 (.A(ALU_OPA[28]),
	.ZN(FE_DBTN13_ALU_OPA_28));
   INV_X1 FE_DBTC12_ALU_OPA_26 (.A(ALU_OPA[26]),
	.ZN(FE_DBTN12_ALU_OPA_26));
   INV_X1 FE_DBTC11_ALU_OPA_24 (.A(FE_OFN117_ALU_OPA_24),
	.ZN(FE_DBTN11_ALU_OPA_24));
   INV_X1 FE_DBTC10_ALU_OPA_22 (.A(ALU_OPA[22]),
	.ZN(FE_DBTN10_ALU_OPA_22));
   INV_X1 FE_DBTC9_ALU_OPA_20 (.A(ALU_OPA[20]),
	.ZN(FE_DBTN9_ALU_OPA_20));
   INV_X1 FE_DBTC8_ALU_OPA_18 (.A(FE_OFN119_ALU_OPA_18),
	.ZN(FE_DBTN8_ALU_OPA_18));
   INV_X1 FE_DBTC7_ALU_OPA_16 (.A(ALU_OPA[16]),
	.ZN(FE_DBTN7_ALU_OPA_16));
   INV_X1 FE_DBTC6_ALU_OPB_3 (.A(ALU_OPB[3]),
	.ZN(FE_DBTN6_ALU_OPB_3));
   INV_X2 FE_DBTC5_ALU_OPB_0 (.A(FE_OFN115_ALU_OPB_0),
	.ZN(FE_DBTN5_ALU_OPB_0));
   INV_X1 FE_DBTC4_n4 (.A(n4),
	.ZN(FE_DBTN4_n4));
   alu_N32_DW01_add_0 add_53 (.A({ ALU_OPA[31],
		FE_OFN116_ALU_OPA_30,
		ALU_OPA[29],
		ALU_OPA[28],
		ALU_OPA[27],
		ALU_OPA[26],
		ALU_OPA[25],
		FE_OFN117_ALU_OPA_24,
		FE_OFN118_ALU_OPA_23,
		ALU_OPA[22],
		ALU_OPA[21],
		ALU_OPA[20],
		ALU_OPA[19],
		FE_OFN119_ALU_OPA_18,
		ALU_OPA[17],
		ALU_OPA[16],
		ALU_OPA[15],
		FE_OFN120_ALU_OPA_14,
		ALU_OPA[13],
		FE_OFN122_ALU_OPA_12,
		ALU_OPA[11],
		FE_OFN121_ALU_OPA_10,
		ALU_OPA[9],
		FE_OFN126_ALU_OPA_8,
		FE_OFN125_ALU_OPA_7,
		FE_OFN127_ALU_OPA_6,
		ALU_OPA[5],
		ALU_OPA[4],
		FE_OFN124_ALU_OPA_3,
		ALU_OPA[2],
		ALU_OPA[1],
		ALU_OPA[0] }),
	.B({ ALU_OPB[31],
		ALU_OPB[30],
		ALU_OPB[29],
		ALU_OPB[28],
		ALU_OPB[27],
		ALU_OPB[26],
		ALU_OPB[25],
		ALU_OPB[24],
		ALU_OPB[23],
		ALU_OPB[22],
		ALU_OPB[21],
		ALU_OPB[20],
		ALU_OPB[19],
		ALU_OPB[18],
		ALU_OPB[17],
		ALU_OPB[16],
		ALU_OPB[15],
		ALU_OPB[14],
		ALU_OPB[13],
		ALU_OPB[12],
		ALU_OPB[11],
		ALU_OPB[10],
		ALU_OPB[9],
		ALU_OPB[8],
		ALU_OPB[7],
		ALU_OPB[6],
		ALU_OPB[5],
		FE_OFN128_ALU_OPB_4,
		ALU_OPB[3],
		ALU_OPB[2],
		ALU_OPB[1],
		FE_OFN115_ALU_OPB_0 }),
	.CI(1'b0),
	.SUM({ N703,
		N702,
		N701,
		N700,
		N699,
		N698,
		N697,
		N696,
		N695,
		N694,
		N693,
		N692,
		N691,
		N690,
		N689,
		N688,
		N687,
		N686,
		N685,
		N684,
		N683,
		N682,
		N681,
		N680,
		N679,
		N678,
		N677,
		N676,
		N675,
		N674,
		N673,
		N672 }));
   alu_N32_DW_cmp_0 lt_47 (.A({ FE_DBTN15_ALU_OPA_31,
		FE_DBTN14_ALU_OPA_30,
		ALU_OPA[29],
		FE_DBTN13_ALU_OPA_28,
		ALU_OPA[27],
		FE_DBTN12_ALU_OPA_26,
		ALU_OPA[25],
		FE_DBTN11_ALU_OPA_24,
		FE_OFN118_ALU_OPA_23,
		FE_DBTN10_ALU_OPA_22,
		ALU_OPA[21],
		FE_DBTN9_ALU_OPA_20,
		ALU_OPA[19],
		FE_DBTN8_ALU_OPA_18,
		ALU_OPA[17],
		FE_DBTN7_ALU_OPA_16,
		ALU_OPA[15],
		FE_OFN120_ALU_OPA_14,
		ALU_OPA[13],
		FE_OFN122_ALU_OPA_12,
		ALU_OPA[11],
		FE_OFN121_ALU_OPA_10,
		ALU_OPA[9],
		FE_OFN126_ALU_OPA_8,
		FE_OFN125_ALU_OPA_7,
		FE_OFN127_ALU_OPA_6,
		FE_OFN123_ALU_OPA_5,
		ALU_OPA[4],
		FE_OFN124_ALU_OPA_3,
		ALU_OPA[2],
		ALU_OPA[1],
		FE_OFN130_ALU_OPA_0 }),
	.B({ ALU_OPB[31],
		ALU_OPB[30],
		ALU_OPB[29],
		ALU_OPB[28],
		ALU_OPB[27],
		ALU_OPB[26],
		ALU_OPB[25],
		ALU_OPB[24],
		ALU_OPB[23],
		ALU_OPB[22],
		ALU_OPB[21],
		ALU_OPB[20],
		ALU_OPB[19],
		ALU_OPB[18],
		ALU_OPB[17],
		ALU_OPB[16],
		ALU_OPB[15],
		ALU_OPB[14],
		ALU_OPB[13],
		ALU_OPB[12],
		ALU_OPB[11],
		ALU_OPB[10],
		ALU_OPB[9],
		ALU_OPB[8],
		ALU_OPB[7],
		ALU_OPB[6],
		ALU_OPB[5],
		FE_OFN128_ALU_OPB_4,
		FE_DBTN6_ALU_OPB_3,
		FE_UNCONNECTED_1,
		ALU_OPB[1],
		FE_OFN115_ALU_OPB_0 }),
	.TC(1'b1),
	.GE_LT(1'b1),
	.GE_GT_EQ(1'b0),
	.GE_LT_GT_LE(N671),
	.n188(n188),
	.n33(ALU_OPB[2]));
   AOI221_X1 U3 (.A(n44),
	.B1(ALU_OPA[2]),
	.B2(n30),
	.C1(FE_OFN124_ALU_OPA_3),
	.C2(n29),
	.ZN(n31));
   AOI221_X1 U5 (.A(n144),
	.B1(ALU_OPA[9]),
	.B2(n91),
	.C1(ALU_OPA[1]),
	.C2(n90),
	.ZN(n58));
   OR3_X1 U11 (.A1(OP[0]),
	.A2(OP[2]),
	.A3(n550),
	.ZN(n4));
   INV_X1 U18 (.A(n304),
	.ZN(n280));
   INV_X1 U19 (.A(n123),
	.ZN(n134));
   NOR2_X1 U20 (.A1(N334),
	.A2(N335),
	.ZN(n317));
   INV_X1 U21 (.A(n83),
	.ZN(n130));
   INV_X1 U25 (.A(n99),
	.ZN(n135));
   XOR2_X1 U28 (.A(n45),
	.B(r422_carry[2]),
	.Z(N332));
   INV_X1 U29 (.A(n110),
	.ZN(n143));
   INV_X1 U30 (.A(n101),
	.ZN(n147));
   INV_X1 U31 (.A(n90),
	.ZN(n129));
   INV_X1 U33 (.A(n91),
	.ZN(n133));
   INV_X1 U34 (.A(n106),
	.ZN(n154));
   INV_X1 U35 (.A(n59),
	.ZN(n146));
   INV_X1 U36 (.A(n121),
	.ZN(n140));
   INV_X2 U37 (.A(n10),
	.ZN(n171));
   INV_X1 U46 (.A(n89),
	.ZN(n149));
   INV_X1 U47 (.A(n47),
	.ZN(n139));
   INV_X1 U48 (.A(n51),
	.ZN(n137));
   INV_X1 U49 (.A(n48),
	.ZN(n138));
   INV_X1 U50 (.A(n84),
	.ZN(n151));
   INV_X1 U51 (.A(n15),
	.ZN(n41));
   INV_X1 U52 (.A(n28),
	.ZN(n44));
   INV_X1 U53 (.A(n22),
	.ZN(n37));
   INV_X1 U54 (.A(n12),
	.ZN(n40));
   INV_X1 U55 (.A(n49),
	.ZN(n153));
   INV_X1 U56 (.A(n54),
	.ZN(n148));
   INV_X1 U57 (.A(n11),
	.ZN(n39));
   INV_X1 U58 (.A(n25),
	.ZN(n38));
   INV_X1 U59 (.A(FE_OFN128_ALU_OPB_4),
	.ZN(n128));
   INV_X1 U60 (.A(ALU_OPA[19]),
	.ZN(n142));
   INV_X1 U61 (.A(ALU_OPA[11]),
	.ZN(n152));
   AND2_X1 U62 (.A1(ALU_OPA[31]),
	.A2(n171),
	.ZN(n9));
   INV_X1 U63 (.A(n46),
	.ZN(n144));
   INV_X1 U64 (.A(n55),
	.ZN(n131));
   INV_X1 U65 (.A(n113),
	.ZN(n141));
   INV_X1 U66 (.A(n16),
	.ZN(n42));
   INV_X1 U67 (.A(n21),
	.ZN(n43));
   INV_X1 U68 (.A(n96),
	.ZN(n145));
   INV_X1 U70 (.A(n52),
	.ZN(n150));
   OR3_X1 U76 (.A1(n550),
	.A2(OP[2]),
	.A3(n549),
	.ZN(n10));
   NOR2_X1 U77 (.A1(n188),
	.A2(FE_OFN115_ALU_OPB_0),
	.ZN(n30));
   NOR2_X1 U78 (.A1(n188),
	.A2(FE_DBTN5_ALU_OPB_0),
	.ZN(n29));
   NOR2_X1 U79 (.A1(FE_OFN115_ALU_OPB_0),
	.A2(ALU_OPB[1]),
	.ZN(n27));
   NOR2_X1 U80 (.A1(FE_DBTN5_ALU_OPB_0),
	.A2(ALU_OPB[1]),
	.ZN(n26));
   AOI22_X1 U81 (.A1(ALU_OPA[28]),
	.A2(n27),
	.B1(ALU_OPA[29]),
	.B2(n26),
	.ZN(n11));
   AOI221_X1 U82 (.A(n39),
	.B1(FE_OFN116_ALU_OPA_30),
	.B2(n30),
	.C1(ALU_OPA[31]),
	.C2(n29),
	.ZN(n14));
   AOI22_X1 U83 (.A1(FE_OFN117_ALU_OPA_24),
	.A2(n27),
	.B1(ALU_OPA[25]),
	.B2(n26),
	.ZN(n12));
   AOI221_X1 U84 (.A(n40),
	.B1(ALU_OPA[26]),
	.B2(n30),
	.C1(ALU_OPA[27]),
	.C2(n29),
	.ZN(n13));
   OAI22_X1 U85 (.A1(n45),
	.A2(n14),
	.B1(ALU_OPB[2]),
	.B2(n13),
	.ZN(n20));
   AOI22_X1 U86 (.A1(ALU_OPA[20]),
	.A2(n27),
	.B1(ALU_OPA[21]),
	.B2(n26),
	.ZN(n15));
   AOI221_X1 U87 (.A(n41),
	.B1(ALU_OPA[22]),
	.B2(n30),
	.C1(FE_OFN118_ALU_OPA_23),
	.C2(n29),
	.ZN(n18));
   AOI22_X1 U88 (.A1(ALU_OPA[16]),
	.A2(n27),
	.B1(ALU_OPA[17]),
	.B2(n26),
	.ZN(n16));
   AOI221_X1 U89 (.A(n42),
	.B1(FE_OFN119_ALU_OPA_18),
	.B2(n30),
	.C1(ALU_OPA[19]),
	.C2(n29),
	.ZN(n17));
   OAI22_X1 U90 (.A1(n18),
	.A2(n45),
	.B1(ALU_OPB[2]),
	.B2(n17),
	.ZN(n19));
   AOI22_X1 U91 (.A1(ALU_OPB[3]),
	.A2(n20),
	.B1(n19),
	.B2(FE_DBTN6_ALU_OPB_3),
	.ZN(n36));
   AOI22_X1 U92 (.A1(FE_OFN122_ALU_OPA_12),
	.A2(n27),
	.B1(ALU_OPA[13]),
	.B2(n26),
	.ZN(n21));
   AOI221_X1 U93 (.A(n43),
	.B1(FE_OFN120_ALU_OPA_14),
	.B2(n30),
	.C1(ALU_OPA[15]),
	.C2(n29),
	.ZN(n24));
   AOI22_X1 U94 (.A1(FE_OFN126_ALU_OPA_8),
	.A2(n27),
	.B1(ALU_OPA[9]),
	.B2(n26),
	.ZN(n22));
   AOI221_X1 U95 (.A(n37),
	.B1(FE_OFN121_ALU_OPA_10),
	.B2(n30),
	.C1(ALU_OPA[11]),
	.C2(n29),
	.ZN(n23));
   OAI22_X1 U96 (.A1(n45),
	.A2(n24),
	.B1(ALU_OPB[2]),
	.B2(n23),
	.ZN(n34));
   AOI22_X1 U97 (.A1(ALU_OPA[4]),
	.A2(n27),
	.B1(FE_OFN123_ALU_OPA_5),
	.B2(n26),
	.ZN(n25));
   AOI221_X1 U98 (.A(n38),
	.B1(FE_OFN127_ALU_OPA_6),
	.B2(n30),
	.C1(FE_OFN125_ALU_OPA_7),
	.C2(n29),
	.ZN(n32));
   AOI22_X1 U99 (.A1(FE_OFN130_ALU_OPA_0),
	.A2(n27),
	.B1(ALU_OPA[1]),
	.B2(n26),
	.ZN(n28));
   OAI22_X1 U100 (.A1(n45),
	.A2(n32),
	.B1(ALU_OPB[2]),
	.B2(n31),
	.ZN(n33));
   AOI22_X1 U101 (.A1(n34),
	.A2(ALU_OPB[3]),
	.B1(n33),
	.B2(FE_DBTN6_ALU_OPB_3),
	.ZN(n35));
   OAI22_X1 U102 (.A1(n36),
	.A2(n128),
	.B1(FE_OFN128_ALU_OPB_4),
	.B2(n35),
	.ZN(N669));
   INV_X2 U103 (.A(ALU_OPB[2]),
	.ZN(n45));
   NAND2_X1 U104 (.A1(n45),
	.A2(FE_DBTN5_ALU_OPB_0),
	.ZN(n103));
   OR2_X1 U105 (.A1(n103),
	.A2(ALU_OPB[1]),
	.ZN(n105));
   NOR2_X1 U106 (.A1(FE_DBTN6_ALU_OPB_3),
	.A2(FE_OFN128_ALU_OPB_4),
	.ZN(n91));
   NOR2_X1 U107 (.A1(ALU_OPB[3]),
	.A2(FE_OFN128_ALU_OPB_4),
	.ZN(n90));
   NOR2_X1 U108 (.A1(n128),
	.A2(ALU_OPB[3]),
	.ZN(n83));
   NAND2_X1 U109 (.A1(FE_OFN128_ALU_OPB_4),
	.A2(ALU_OPB[3]),
	.ZN(n55));
   AOI22_X1 U110 (.A1(ALU_OPA[17]),
	.A2(n83),
	.B1(ALU_OPA[25]),
	.B2(n131),
	.ZN(n46));
   NOR2_X1 U111 (.A1(n45),
	.A2(FE_OFN115_ALU_OPB_0),
	.ZN(n123));
   OAI22_X1 U112 (.A1(n55),
	.A2(ALU_OPA[29]),
	.B1(n130),
	.B2(ALU_OPA[21]),
	.ZN(n47));
   OAI221_X1 U113 (.A(n139),
	.B1(ALU_OPA[13]),
	.B2(n133),
	.C1(FE_OFN123_ALU_OPA_5),
	.C2(n129),
	.ZN(n59));
   OAI22_X1 U114 (.A1(n55),
	.A2(FE_OFN116_ALU_OPA_30),
	.B1(n130),
	.B2(ALU_OPA[22]),
	.ZN(n48));
   OAI221_X1 U115 (.A(n138),
	.B1(FE_OFN120_ALU_OPA_14),
	.B2(n133),
	.C1(FE_OFN127_ALU_OPA_6),
	.C2(n129),
	.ZN(n64));
   OAI22_X1 U116 (.A1(ALU_OPA[2]),
	.A2(n129),
	.B1(FE_OFN121_ALU_OPA_10),
	.B2(n133),
	.ZN(n49));
   OAI221_X1 U117 (.A(n153),
	.B1(n55),
	.B2(ALU_OPA[26]),
	.C1(n130),
	.C2(FE_OFN119_ALU_OPA_18),
	.ZN(n50));
   AOI22_X1 U118 (.A1(ALU_OPB[2]),
	.A2(n64),
	.B1(n45),
	.B2(n50),
	.ZN(n61));
   AOI22_X1 U119 (.A1(n123),
	.A2(n146),
	.B1(FE_OFN115_ALU_OPB_0),
	.B2(n61),
	.ZN(n57));
   OAI22_X1 U120 (.A1(n55),
	.A2(ALU_OPA[31]),
	.B1(n130),
	.B2(FE_OFN118_ALU_OPA_23),
	.ZN(n51));
   OAI221_X1 U121 (.A(n137),
	.B1(ALU_OPA[15]),
	.B2(n133),
	.C1(FE_OFN125_ALU_OPA_7),
	.C2(n129),
	.ZN(n67));
   AOI22_X1 U122 (.A1(n352),
	.A2(ALU_OPB[3]),
	.B1(n142),
	.B2(FE_DBTN6_ALU_OPB_3),
	.ZN(n116));
   OAI22_X1 U123 (.A1(FE_OFN124_ALU_OPA_3),
	.A2(n129),
	.B1(ALU_OPA[11]),
	.B2(n133),
	.ZN(n52));
   OAI21_X1 U124 (.A(n150),
	.B1(n116),
	.B2(n128),
	.ZN(n53));
   AOI22_X1 U125 (.A1(ALU_OPB[2]),
	.A2(n67),
	.B1(n45),
	.B2(n53),
	.ZN(n62));
   OAI222_X1 U126 (.A1(FE_OFN126_ALU_OPA_8),
	.A2(n129),
	.B1(FE_OFN117_ALU_OPA_24),
	.B2(n130),
	.C1(ALU_OPA[16]),
	.C2(FE_DBTN6_ALU_OPB_3),
	.ZN(n71));
   OAI22_X1 U127 (.A1(ALU_OPA[4]),
	.A2(n129),
	.B1(FE_OFN122_ALU_OPA_12),
	.B2(n133),
	.ZN(n54));
   OAI221_X1 U128 (.A(n148),
	.B1(n55),
	.B2(ALU_OPA[28]),
	.C1(n130),
	.C2(ALU_OPA[20]),
	.ZN(n56));
   AOI22_X1 U129 (.A1(ALU_OPB[2]),
	.A2(n71),
	.B1(n45),
	.B2(n56),
	.ZN(n60));
   AOI22_X1 U130 (.A1(FE_DBTN5_ALU_OPB_0),
	.A2(n62),
	.B1(n60),
	.B2(FE_OFN115_ALU_OPB_0),
	.ZN(n66));
   OAI222_X1 U131 (.A1(n105),
	.A2(n58),
	.B1(ALU_OPB[1]),
	.B2(n57),
	.C1(n188),
	.C2(n66),
	.ZN(N665));
   OAI222_X1 U132 (.A1(ALU_OPA[9]),
	.A2(n129),
	.B1(ALU_OPA[25]),
	.B2(n130),
	.C1(ALU_OPA[17]),
	.C2(FE_DBTN6_ALU_OPB_3),
	.ZN(n75));
   AOI22_X1 U133 (.A1(n45),
	.A2(n59),
	.B1(ALU_OPB[2]),
	.B2(n75),
	.ZN(n65));
   OAI22_X1 U134 (.A1(FE_OFN115_ALU_OPB_0),
	.A2(n60),
	.B1(FE_DBTN5_ALU_OPB_0),
	.B2(n65),
	.ZN(n69));
   AOI22_X1 U135 (.A1(FE_OFN115_ALU_OPB_0),
	.A2(n62),
	.B1(n61),
	.B2(FE_DBTN5_ALU_OPB_0),
	.ZN(n63));
   OAI22_X1 U136 (.A1(n69),
	.A2(n188),
	.B1(ALU_OPB[1]),
	.B2(n63),
	.ZN(N661));
   OAI222_X1 U137 (.A1(FE_OFN121_ALU_OPA_10),
	.A2(n129),
	.B1(ALU_OPA[26]),
	.B2(n130),
	.C1(FE_OFN119_ALU_OPA_18),
	.C2(FE_DBTN6_ALU_OPB_3),
	.ZN(n79));
   AOI22_X1 U138 (.A1(n45),
	.A2(n64),
	.B1(ALU_OPB[2]),
	.B2(n79),
	.ZN(n68));
   OAI22_X1 U139 (.A1(FE_OFN115_ALU_OPB_0),
	.A2(n65),
	.B1(FE_DBTN5_ALU_OPB_0),
	.B2(n68),
	.ZN(n73));
   OAI22_X1 U140 (.A1(n73),
	.A2(n188),
	.B1(ALU_OPB[1]),
	.B2(n66),
	.ZN(N657));
   OAI222_X1 U141 (.A1(ALU_OPA[11]),
	.A2(n129),
	.B1(ALU_OPA[27]),
	.B2(n130),
	.C1(ALU_OPA[19]),
	.C2(FE_DBTN6_ALU_OPB_3),
	.ZN(n84));
   AOI22_X1 U142 (.A1(n45),
	.A2(n67),
	.B1(ALU_OPB[2]),
	.B2(n84),
	.ZN(n72));
   OAI22_X1 U143 (.A1(FE_OFN115_ALU_OPB_0),
	.A2(n68),
	.B1(FE_DBTN5_ALU_OPB_0),
	.B2(n72),
	.ZN(n77));
   OAI22_X1 U144 (.A1(ALU_OPB[1]),
	.A2(n69),
	.B1(n77),
	.B2(n188),
	.ZN(N653));
   OAI222_X1 U145 (.A1(FE_DBTN6_ALU_OPB_3),
	.A2(ALU_OPA[20]),
	.B1(n130),
	.B2(ALU_OPA[28]),
	.C1(n129),
	.C2(FE_OFN122_ALU_OPA_12),
	.ZN(n70));
   AOI22_X1 U146 (.A1(n45),
	.A2(n71),
	.B1(ALU_OPB[2]),
	.B2(n70),
	.ZN(n76));
   OAI22_X1 U147 (.A1(FE_DBTN5_ALU_OPB_0),
	.A2(n76),
	.B1(FE_OFN115_ALU_OPB_0),
	.B2(n72),
	.ZN(n82));
   OAI22_X1 U148 (.A1(ALU_OPB[1]),
	.A2(n73),
	.B1(n82),
	.B2(n188),
	.ZN(N649));
   OAI222_X1 U149 (.A1(FE_DBTN6_ALU_OPB_3),
	.A2(ALU_OPA[21]),
	.B1(n130),
	.B2(ALU_OPA[29]),
	.C1(n129),
	.C2(ALU_OPA[13]),
	.ZN(n74));
   AOI22_X1 U150 (.A1(n45),
	.A2(n75),
	.B1(ALU_OPB[2]),
	.B2(n74),
	.ZN(n80));
   AOI22_X1 U151 (.A1(FE_DBTN5_ALU_OPB_0),
	.A2(n76),
	.B1(n80),
	.B2(FE_OFN115_ALU_OPB_0),
	.ZN(n86));
   OAI22_X1 U152 (.A1(ALU_OPB[1]),
	.A2(n77),
	.B1(n188),
	.B2(n86),
	.ZN(N645));
   OAI222_X1 U153 (.A1(FE_DBTN6_ALU_OPB_3),
	.A2(ALU_OPA[22]),
	.B1(n130),
	.B2(FE_OFN116_ALU_OPA_30),
	.C1(n129),
	.C2(FE_OFN120_ALU_OPA_14),
	.ZN(n78));
   AOI22_X1 U154 (.A1(n45),
	.A2(n79),
	.B1(ALU_OPB[2]),
	.B2(n78),
	.ZN(n85));
   AOI22_X1 U155 (.A1(FE_OFN115_ALU_OPB_0),
	.A2(n85),
	.B1(n80),
	.B2(FE_DBTN5_ALU_OPB_0),
	.ZN(n81));
   OAI22_X1 U156 (.A1(ALU_OPB[1]),
	.A2(n82),
	.B1(n188),
	.B2(n81),
	.ZN(N641));
   NAND2_X1 U157 (.A1(ALU_OPB[2]),
	.A2(FE_OFN115_ALU_OPB_0),
	.ZN(n115));
   OR2_X1 U158 (.A1(n188),
	.A2(n115),
	.ZN(n125));
   AOI222_X1 U159 (.A1(FE_OFN118_ALU_OPA_23),
	.A2(ALU_OPB[3]),
	.B1(ALU_OPA[31]),
	.B2(n83),
	.C1(ALU_OPA[15]),
	.C2(n90),
	.ZN(n88));
   NOR2_X1 U160 (.A1(FE_DBTN5_ALU_OPB_0),
	.A2(ALU_OPB[2]),
	.ZN(n99));
   AOI22_X1 U161 (.A1(n99),
	.A2(n151),
	.B1(n85),
	.B2(FE_DBTN5_ALU_OPB_0),
	.ZN(n87));
   OAI222_X1 U162 (.A1(n125),
	.A2(n88),
	.B1(n188),
	.B2(n87),
	.C1(ALU_OPB[1]),
	.C2(n86),
	.ZN(N637));
   AOI222_X1 U163 (.A1(ALU_OPA[25]),
	.A2(FE_OFN128_ALU_OPB_4),
	.B1(ALU_OPA[17]),
	.B2(n91),
	.C1(ALU_OPA[9]),
	.C2(n90),
	.ZN(n95));
   AOI222_X1 U164 (.A1(n90),
	.A2(FE_OFN121_ALU_OPA_10),
	.B1(n91),
	.B2(FE_OFN119_ALU_OPA_18),
	.C1(FE_OFN128_ALU_OPB_4),
	.C2(ALU_OPA[26]),
	.ZN(n106));
   OAI222_X1 U165 (.A1(ALU_OPA[13]),
	.A2(n129),
	.B1(ALU_OPA[21]),
	.B2(n133),
	.C1(ALU_OPA[29]),
	.C2(n128),
	.ZN(n101));
   OAI222_X1 U166 (.A1(FE_OFN120_ALU_OPA_14),
	.A2(n129),
	.B1(ALU_OPA[22]),
	.B2(n133),
	.C1(FE_OFN116_ALU_OPA_30),
	.C2(n128),
	.ZN(n98));
   AOI22_X1 U167 (.A1(FE_DBTN5_ALU_OPB_0),
	.A2(n101),
	.B1(FE_OFN115_ALU_OPB_0),
	.B2(n98),
	.ZN(n108));
   AOI22_X1 U168 (.A1(n154),
	.A2(n99),
	.B1(ALU_OPB[2]),
	.B2(n108),
	.ZN(n94));
   OAI222_X1 U169 (.A1(FE_OFN122_ALU_OPA_12),
	.A2(n129),
	.B1(ALU_OPA[20]),
	.B2(n133),
	.C1(ALU_OPA[28]),
	.C2(n128),
	.ZN(n89));
   AOI222_X1 U170 (.A1(FE_OFN128_ALU_OPB_4),
	.A2(n352),
	.B1(n91),
	.B2(n142),
	.C1(n90),
	.C2(n152),
	.ZN(n93));
   OAI22_X1 U171 (.A1(ALU_OPA[15]),
	.A2(n129),
	.B1(FE_OFN118_ALU_OPA_23),
	.B2(n133),
	.ZN(n96));
   OAI22_X1 U172 (.A1(n133),
	.A2(FE_OFN117_ALU_OPA_24),
	.B1(n129),
	.B2(ALU_OPA[16]),
	.ZN(n92));
   AOI222_X1 U173 (.A1(FE_DBTN5_ALU_OPB_0),
	.A2(n96),
	.B1(n92),
	.B2(FE_OFN115_ALU_OPB_0),
	.C1(FE_DBTN15_ALU_OPA_31),
	.C2(FE_OFN128_ALU_OPB_4),
	.ZN(n114));
   OAI222_X1 U174 (.A1(n149),
	.A2(n135),
	.B1(n103),
	.B2(n93),
	.C1(n114),
	.C2(n45),
	.ZN(n109));
   OAI222_X1 U175 (.A1(n105),
	.A2(n95),
	.B1(ALU_OPB[1]),
	.B2(n94),
	.C1(n109),
	.C2(n188),
	.ZN(N633));
   OAI222_X1 U176 (.A1(n129),
	.A2(n152),
	.B1(n133),
	.B2(n142),
	.C1(n128),
	.C2(n352),
	.ZN(n100));
   OAI21_X1 U177 (.A(n145),
	.B1(n128),
	.B2(ALU_OPA[31]),
	.ZN(n97));
   AOI22_X1 U178 (.A1(FE_DBTN5_ALU_OPB_0),
	.A2(n98),
	.B1(FE_OFN115_ALU_OPB_0),
	.B2(n97),
	.ZN(n111));
   AOI22_X1 U179 (.A1(n100),
	.A2(n99),
	.B1(ALU_OPB[2]),
	.B2(n111),
	.ZN(n104));
   OAI22_X1 U180 (.A1(ALU_OPA[25]),
	.A2(FE_DBTN6_ALU_OPB_3),
	.B1(ALU_OPA[17]),
	.B2(ALU_OPB[3]),
	.ZN(n107));
   OAI22_X1 U181 (.A1(ALU_OPB[3]),
	.A2(ALU_OPA[16]),
	.B1(FE_DBTN6_ALU_OPB_3),
	.B2(FE_OFN117_ALU_OPA_24),
	.ZN(n102));
   AOI22_X1 U182 (.A1(FE_OFN115_ALU_OPB_0),
	.A2(n107),
	.B1(FE_DBTN5_ALU_OPB_0),
	.B2(n102),
	.ZN(n118));
   OAI222_X1 U183 (.A1(n147),
	.A2(n135),
	.B1(n149),
	.B2(n103),
	.C1(n45),
	.C2(n118),
	.ZN(n112));
   OAI222_X1 U184 (.A1(n106),
	.A2(n105),
	.B1(ALU_OPB[1]),
	.B2(n104),
	.C1(n112),
	.C2(n188),
	.ZN(N629));
   OAI22_X1 U185 (.A1(ALU_OPA[26]),
	.A2(FE_DBTN6_ALU_OPB_3),
	.B1(FE_OFN119_ALU_OPA_18),
	.B2(ALU_OPB[3]),
	.ZN(n110));
   AOI22_X1 U186 (.A1(FE_DBTN5_ALU_OPB_0),
	.A2(n107),
	.B1(FE_OFN115_ALU_OPB_0),
	.B2(n110),
	.ZN(n122));
   AOI22_X1 U187 (.A1(n45),
	.A2(n108),
	.B1(n122),
	.B2(ALU_OPB[2]),
	.ZN(n117));
   OAI22_X1 U188 (.A1(ALU_OPB[1]),
	.A2(n109),
	.B1(n188),
	.B2(n117),
	.ZN(N625));
   OAI222_X1 U189 (.A1(n134),
	.A2(n143),
	.B1(n116),
	.B2(n115),
	.C1(ALU_OPB[2]),
	.C2(n111),
	.ZN(n119));
   OAI22_X1 U190 (.A1(ALU_OPB[1]),
	.A2(n112),
	.B1(n119),
	.B2(n188),
	.ZN(N621));
   OAI22_X1 U191 (.A1(ALU_OPA[28]),
	.A2(FE_DBTN6_ALU_OPB_3),
	.B1(ALU_OPA[20]),
	.B2(ALU_OPB[3]),
	.ZN(n113));
   OAI222_X1 U192 (.A1(n116),
	.A2(n134),
	.B1(n141),
	.B2(n115),
	.C1(ALU_OPB[2]),
	.C2(n114),
	.ZN(n124));
   OAI22_X1 U193 (.A1(n124),
	.A2(n188),
	.B1(ALU_OPB[1]),
	.B2(n117),
	.ZN(N617));
   AOI22_X1 U194 (.A1(ALU_OPB[3]),
	.A2(ALU_OPA[29]),
	.B1(FE_DBTN6_ALU_OPB_3),
	.B2(ALU_OPA[21]),
	.ZN(n121));
   AOI22_X1 U195 (.A1(n123),
	.A2(n141),
	.B1(n118),
	.B2(n45),
	.ZN(n120));
   OAI222_X1 U196 (.A1(n121),
	.A2(n125),
	.B1(n188),
	.B2(n120),
	.C1(ALU_OPB[1]),
	.C2(n119),
	.ZN(N613));
   AOI22_X1 U197 (.A1(n140),
	.A2(n123),
	.B1(n122),
	.B2(n45),
	.ZN(n127));
   AOI22_X1 U198 (.A1(ALU_OPA[22]),
	.A2(FE_DBTN6_ALU_OPB_3),
	.B1(FE_OFN116_ALU_OPA_30),
	.B2(ALU_OPB[3]),
	.ZN(n126));
   OAI222_X1 U199 (.A1(n188),
	.A2(n127),
	.B1(n126),
	.B2(n125),
	.C1(ALU_OPB[1]),
	.C2(n124),
	.ZN(N591));
   INV_X1 U211 (.A(n9),
	.ZN(n170));
   INV_X1 U212 (.A(ALU_OPB[1]),
	.ZN(n188));
   AND2_X1 U213 (.A1(r422_carry[4]),
	.A2(n128),
	.ZN(N335));
   XOR2_X1 U214 (.A(n128),
	.B(r422_carry[4]),
	.Z(N334));
   AND2_X1 U215 (.A1(r422_carry[3]),
	.A2(FE_DBTN6_ALU_OPB_3),
	.ZN(r422_carry[4]));
   XOR2_X1 U216 (.A(FE_DBTN6_ALU_OPB_3),
	.B(r422_carry[3]),
	.Z(N333));
   AND2_X1 U217 (.A1(r422_carry[2]),
	.A2(n45),
	.ZN(r422_carry[3]));
   AND2_X1 U218 (.A1(FE_DBTN5_ALU_OPB_0),
	.A2(n188),
	.ZN(r422_carry[2]));
   XOR2_X1 U219 (.A(n188),
	.B(FE_DBTN5_ALU_OPB_0),
	.Z(N331));
   NAND3_X1 U220 (.A1(n189),
	.A2(n190),
	.A3(n191),
	.ZN(ALU_OUT[9]));
   MUX2_X1 U221 (.A(n192),
	.B(n170),
	.S(n193),
	.Z(n191));
   AOI21_X1 U222 (.A(n194),
	.B1(N331),
	.B2(N333),
	.ZN(n193));
   NAND2_X1 U223 (.A1(N633),
	.A2(n171),
	.ZN(n192));
   NAND2_X1 U224 (.A1(N681),
	.A2(FE_OFN34_n198),
	.ZN(n190));
   MUX2_X1 U225 (.A(n199),
	.B(n200),
	.S(ALU_OPB[9]),
	.Z(n189));
   MUX2_X1 U226 (.A(n4),
	.B(n201),
	.S(ALU_OPA[9]),
	.Z(n200));
   NAND2_X1 U227 (.A1(ALU_OPA[9]),
	.A2(FE_OFN42_FE_DBTN4_n4),
	.ZN(n199));
   NAND3_X1 U228 (.A1(n202),
	.A2(n203),
	.A3(n204),
	.ZN(ALU_OUT[8]));
   MUX2_X1 U229 (.A(n170),
	.B(n205),
	.S(n206),
	.Z(n204));
   NOR2_X1 U230 (.A1(n207),
	.A2(n208),
	.ZN(n206));
   NOR3_X1 U231 (.A1(n209),
	.A2(N332),
	.A3(n210),
	.ZN(n207));
   NAND2_X1 U232 (.A1(N637),
	.A2(n171),
	.ZN(n205));
   NAND2_X1 U233 (.A1(N680),
	.A2(FE_OFN34_n198),
	.ZN(n203));
   MUX2_X1 U234 (.A(n211),
	.B(n212),
	.S(ALU_OPB[8]),
	.Z(n202));
   MUX2_X1 U235 (.A(n4),
	.B(n201),
	.S(FE_OFN126_ALU_OPA_8),
	.Z(n212));
   NAND2_X1 U236 (.A1(FE_OFN126_ALU_OPA_8),
	.A2(FE_OFN42_FE_DBTN4_n4),
	.ZN(n211));
   NAND3_X1 U237 (.A1(n213),
	.A2(n214),
	.A3(n215),
	.ZN(ALU_OUT[7]));
   MUX2_X1 U238 (.A(n216),
	.B(n170),
	.S(n208),
	.Z(n215));
   NAND2_X1 U239 (.A1(N641),
	.A2(n171),
	.ZN(n216));
   NAND2_X1 U240 (.A1(N679),
	.A2(FE_OFN34_n198),
	.ZN(n214));
   MUX2_X1 U241 (.A(n217),
	.B(n218),
	.S(ALU_OPB[7]),
	.Z(n213));
   MUX2_X1 U242 (.A(n4),
	.B(n201),
	.S(FE_OFN125_ALU_OPA_7),
	.Z(n218));
   NAND2_X1 U243 (.A1(FE_OFN125_ALU_OPA_7),
	.A2(FE_OFN42_FE_DBTN4_n4),
	.ZN(n217));
   NAND3_X1 U244 (.A1(n219),
	.A2(n220),
	.A3(n221),
	.ZN(ALU_OUT[6]));
   MUX2_X1 U245 (.A(n222),
	.B(n170),
	.S(n223),
	.Z(n221));
   OAI21_X1 U246 (.A(n225),
	.B1(n224),
	.B2(FE_OFN115_ALU_OPB_0),
	.ZN(n223));
   NAND2_X1 U247 (.A1(N645),
	.A2(n171),
	.ZN(n222));
   NAND2_X1 U248 (.A1(N678),
	.A2(FE_OFN34_n198),
	.ZN(n220));
   MUX2_X1 U249 (.A(n226),
	.B(n227),
	.S(ALU_OPB[6]),
	.Z(n219));
   MUX2_X1 U250 (.A(n4),
	.B(n201),
	.S(FE_OFN127_ALU_OPA_6),
	.Z(n227));
   NAND2_X1 U251 (.A1(FE_OFN127_ALU_OPA_6),
	.A2(FE_OFN42_FE_DBTN4_n4),
	.ZN(n226));
   NAND3_X1 U252 (.A1(n228),
	.A2(n229),
	.A3(n230),
	.ZN(ALU_OUT[5]));
   MUX2_X1 U253 (.A(n170),
	.B(n231),
	.S(n225),
	.Z(n230));
   AOI21_X1 U254 (.A(n233),
	.B1(n232),
	.B2(n208),
	.ZN(n225));
   NAND2_X1 U255 (.A1(N649),
	.A2(n171),
	.ZN(n231));
   NAND2_X1 U256 (.A1(N677),
	.A2(FE_OFN34_n198),
	.ZN(n229));
   MUX2_X1 U257 (.A(n234),
	.B(n235),
	.S(ALU_OPB[5]),
	.Z(n228));
   MUX2_X1 U258 (.A(n4),
	.B(n201),
	.S(ALU_OPA[5]),
	.Z(n235));
   NAND2_X1 U259 (.A1(ALU_OPA[5]),
	.A2(FE_OFN42_FE_DBTN4_n4),
	.ZN(n234));
   NAND3_X1 U260 (.A1(n236),
	.A2(n237),
	.A3(n238),
	.ZN(ALU_OUT[4]));
   MUX2_X1 U261 (.A(n170),
	.B(n239),
	.S(n240),
	.Z(n238));
   AOI21_X1 U262 (.A(n233),
	.B1(n208),
	.B2(n241),
	.ZN(n240));
   INV_X1 U263 (.A(n224),
	.ZN(n208));
   NAND2_X1 U264 (.A1(N653),
	.A2(n171),
	.ZN(n239));
   NAND2_X1 U265 (.A1(N676),
	.A2(FE_OFN34_n198),
	.ZN(n237));
   MUX2_X1 U266 (.A(n242),
	.B(n243),
	.S(ALU_OPB[4]),
	.Z(n236));
   MUX2_X1 U267 (.A(n4),
	.B(n201),
	.S(ALU_OPA[4]),
	.Z(n243));
   NAND2_X1 U268 (.A1(ALU_OPA[4]),
	.A2(FE_OFN42_FE_DBTN4_n4),
	.ZN(n242));
   NAND3_X1 U269 (.A1(n244),
	.A2(n245),
	.A3(n246),
	.ZN(ALU_OUT[3]));
   MUX2_X1 U270 (.A(n247),
	.B(n170),
	.S(n233),
	.Z(n246));
   NAND2_X1 U271 (.A1(N657),
	.A2(n171),
	.ZN(n247));
   NAND2_X1 U272 (.A1(N675),
	.A2(FE_OFN34_n198),
	.ZN(n245));
   MUX2_X1 U273 (.A(n248),
	.B(n249),
	.S(ALU_OPB[3]),
	.Z(n244));
   MUX2_X1 U274 (.A(n4),
	.B(n201),
	.S(FE_OFN124_ALU_OPA_3),
	.Z(n249));
   NAND2_X1 U275 (.A1(FE_OFN124_ALU_OPA_3),
	.A2(FE_OFN42_FE_DBTN4_n4),
	.ZN(n248));
   NAND2_X1 U276 (.A1(n250),
	.A2(n251),
	.ZN(ALU_OUT[31]));
   MUX2_X1 U277 (.A(n252),
	.B(n253),
	.S(ALU_OPB[31]),
	.Z(n251));
   MUX2_X1 U278 (.A(n4),
	.B(n201),
	.S(ALU_OPA[31]),
	.Z(n253));
   NAND2_X1 U279 (.A1(ALU_OPA[31]),
	.A2(FE_DBTN4_n4),
	.ZN(n252));
   AOI21_X1 U280 (.A(n9),
	.B1(N703),
	.B2(FE_OFN34_n198),
	.ZN(n250));
   INV_X1 U281 (.A(n254),
	.ZN(ALU_OUT[30]));
   AOI221_X1 U282 (.A(n256),
	.B1(n9),
	.B2(n255),
	.C1(N702),
	.C2(FE_OFN34_n198),
	.ZN(n254));
   MUX2_X1 U283 (.A(n257),
	.B(n258),
	.S(FE_OFN116_ALU_OPA_30),
	.Z(n256));
   OAI21_X1 U284 (.A(n259),
	.B1(n10),
	.B2(n255),
	.ZN(n258));
   MUX2_X1 U285 (.A(n4),
	.B(n201),
	.S(ALU_OPB[30]),
	.Z(n259));
   AND2_X1 U286 (.A1(FE_DBTN4_n4),
	.A2(ALU_OPB[30]),
	.ZN(n257));
   NAND2_X1 U287 (.A1(n260),
	.A2(FE_DBTN5_ALU_OPB_0),
	.ZN(n255));
   NAND2_X1 U288 (.A1(n261),
	.A2(n262),
	.ZN(n260));
   NAND3_X1 U289 (.A1(n263),
	.A2(N332),
	.A3(N334),
	.ZN(n262));
   NAND3_X1 U290 (.A1(n264),
	.A2(n265),
	.A3(n266),
	.ZN(ALU_OUT[2]));
   MUX2_X1 U291 (.A(n170),
	.B(n267),
	.S(n268),
	.Z(n266));
   OAI21_X1 U292 (.A(n233),
	.B1(FE_DBTN5_ALU_OPB_0),
	.B2(n232),
	.ZN(n268));
   NAND2_X1 U293 (.A1(N661),
	.A2(n171),
	.ZN(n267));
   NAND2_X1 U294 (.A1(N674),
	.A2(FE_OFN34_n198),
	.ZN(n265));
   MUX2_X1 U295 (.A(n269),
	.B(n270),
	.S(ALU_OPB[2]),
	.Z(n264));
   MUX2_X1 U296 (.A(n4),
	.B(n201),
	.S(ALU_OPA[2]),
	.Z(n270));
   NAND2_X1 U297 (.A1(ALU_OPA[2]),
	.A2(FE_OFN42_FE_DBTN4_n4),
	.ZN(n269));
   OAI221_X1 U298 (.A(n273),
	.B1(n10),
	.B2(n271),
	.C1(n272),
	.C2(n170),
	.ZN(ALU_OUT[29]));
   AOI21_X1 U299 (.A(n274),
	.B1(N701),
	.B2(FE_OFN34_n198),
	.ZN(n273));
   MUX2_X1 U300 (.A(n275),
	.B(n276),
	.S(ALU_OPB[29]),
	.Z(n274));
   MUX2_X1 U301 (.A(FE_OFN42_FE_DBTN4_n4),
	.B(n277),
	.S(ALU_OPA[29]),
	.Z(n276));
   NOR2_X1 U302 (.A1(n4),
	.A2(n278),
	.ZN(n275));
   AOI211_X1 U303 (.A(n279),
	.B(n280),
	.C1(n232),
	.C2(n261),
	.ZN(n272));
   NAND2_X1 U304 (.A1(n281),
	.A2(n282),
	.ZN(n271));
   OAI21_X1 U305 (.A(n261),
	.B1(n283),
	.B2(n284),
	.ZN(n281));
   NAND4_X1 U306 (.A1(n285),
	.A2(n286),
	.A3(n287),
	.A4(n288),
	.ZN(ALU_OUT[28]));
   OR3_X1 U307 (.A1(n10),
	.A2(n289),
	.A3(n290),
	.ZN(n288));
   OAI21_X1 U308 (.A(n9),
	.B1(n291),
	.B2(n290),
	.ZN(n287));
   NAND2_X1 U309 (.A1(n292),
	.A2(n210),
	.ZN(n290));
   OAI21_X1 U310 (.A(n261),
	.B1(n241),
	.B2(n283),
	.ZN(n292));
   NAND2_X1 U311 (.A1(N700),
	.A2(FE_OFN34_n198),
	.ZN(n286));
   MUX2_X1 U312 (.A(n293),
	.B(n294),
	.S(ALU_OPB[28]),
	.Z(n285));
   MUX2_X1 U313 (.A(n4),
	.B(n201),
	.S(ALU_OPA[28]),
	.Z(n294));
   NAND2_X1 U314 (.A1(ALU_OPA[28]),
	.A2(FE_DBTN4_n4),
	.ZN(n293));
   NAND3_X1 U315 (.A1(n295),
	.A2(n296),
	.A3(n297),
	.ZN(ALU_OUT[27]));
   AOI221_X1 U316 (.A(n300),
	.B1(n9),
	.B2(n279),
	.C1(n298),
	.C2(n299),
	.ZN(n297));
   NOR4_X1 U317 (.A1(ALU_OPB[2]),
	.A2(n301),
	.A3(n302),
	.A4(n10),
	.ZN(n300));
   AOI221_X1 U318 (.A(n303),
	.B1(n291),
	.B2(FE_OFN116_ALU_OPA_30),
	.C1(ALU_OPA[27]),
	.C2(n299),
	.ZN(n301));
   OAI22_X1 U319 (.A1(n278),
	.A2(n304),
	.B1(n305),
	.B2(FE_DBTN13_ALU_OPA_28),
	.ZN(n303));
   OAI21_X1 U320 (.A(n307),
	.B1(N335),
	.B2(N332),
	.ZN(n279));
   NAND2_X1 U321 (.A1(N699),
	.A2(FE_OFN34_n198),
	.ZN(n296));
   MUX2_X1 U322 (.A(n308),
	.B(n309),
	.S(ALU_OPB[27]),
	.Z(n295));
   MUX2_X1 U323 (.A(n4),
	.B(n201),
	.S(ALU_OPA[27]),
	.Z(n309));
   NAND2_X1 U324 (.A1(ALU_OPA[27]),
	.A2(FE_DBTN4_n4),
	.ZN(n308));
   NAND3_X1 U325 (.A1(n310),
	.A2(n311),
	.A3(n312),
	.ZN(ALU_OUT[26]));
   AOI22_X1 U326 (.A1(n298),
	.A2(n313),
	.B1(N698),
	.B2(FE_OFN34_n198),
	.ZN(n312));
   MUX2_X1 U327 (.A(n170),
	.B(n314),
	.S(n315),
	.Z(n311));
   AOI21_X1 U328 (.A(n317),
	.B1(n316),
	.B2(n283),
	.ZN(n315));
   NOR2_X1 U329 (.A1(N335),
	.A2(n263),
	.ZN(n316));
   NAND2_X1 U330 (.A1(n171),
	.A2(n318),
	.ZN(n314));
   OAI22_X1 U331 (.A1(n319),
	.A2(n320),
	.B1(ALU_OPB[2]),
	.B2(n321),
	.ZN(n318));
   AOI222_X1 U332 (.A1(n291),
	.A2(ALU_OPA[29]),
	.B1(ALU_OPA[27]),
	.B2(n313),
	.C1(n280),
	.C2(ALU_OPA[28]),
	.ZN(n321));
   MUX2_X1 U333 (.A(n322),
	.B(n323),
	.S(ALU_OPB[26]),
	.Z(n310));
   MUX2_X1 U334 (.A(n4),
	.B(n201),
	.S(ALU_OPA[26]),
	.Z(n323));
   NAND2_X1 U335 (.A1(ALU_OPA[26]),
	.A2(FE_DBTN4_n4),
	.ZN(n322));
   NAND3_X1 U336 (.A1(n324),
	.A2(n325),
	.A3(n326),
	.ZN(ALU_OUT[25]));
   AOI22_X1 U337 (.A1(n298),
	.A2(n280),
	.B1(N697),
	.B2(FE_OFN34_n198),
	.ZN(n326));
   MUX2_X1 U338 (.A(n170),
	.B(n327),
	.S(n328),
	.Z(n325));
   OAI21_X1 U339 (.A(n302),
	.B1(n284),
	.B2(n329),
	.ZN(n328));
   AOI21_X1 U340 (.A(N335),
	.B1(N334),
	.B2(n330),
	.ZN(n302));
   NAND2_X1 U341 (.A1(n171),
	.A2(n331),
	.ZN(n327));
   OAI222_X1 U342 (.A1(n332),
	.A2(n320),
	.B1(ALU_OPB[2]),
	.B2(n333),
	.C1(n319),
	.C2(n305),
	.ZN(n331));
   AOI22_X1 U343 (.A1(ALU_OPA[27]),
	.A2(n280),
	.B1(n291),
	.B2(ALU_OPA[28]),
	.ZN(n333));
   MUX2_X1 U344 (.A(n334),
	.B(n335),
	.S(ALU_OPB[25]),
	.Z(n324));
   MUX2_X1 U345 (.A(n4),
	.B(n201),
	.S(ALU_OPA[25]),
	.Z(n335));
   NAND2_X1 U346 (.A1(ALU_OPA[25]),
	.A2(FE_DBTN4_n4),
	.ZN(n334));
   NAND2_X1 U347 (.A1(n336),
	.A2(n337),
	.ZN(ALU_OUT[24]));
   MUX2_X1 U348 (.A(n338),
	.B(n339),
	.S(ALU_OPB[24]),
	.Z(n337));
   MUX2_X1 U349 (.A(n4),
	.B(n201),
	.S(FE_OFN117_ALU_OPA_24),
	.Z(n339));
   NAND2_X1 U350 (.A1(FE_OFN117_ALU_OPA_24),
	.A2(FE_DBTN4_n4),
	.ZN(n338));
   AOI21_X1 U351 (.A(n340),
	.B1(N696),
	.B2(FE_OFN34_n198),
	.ZN(n336));
   MUX2_X1 U352 (.A(n9),
	.B(n341),
	.S(n342),
	.Z(n340));
   NOR2_X1 U353 (.A1(n343),
	.A2(n344),
	.ZN(n342));
   NOR3_X1 U354 (.A1(n209),
	.A2(N335),
	.A3(N332),
	.ZN(n343));
   INV_X1 U355 (.A(n345),
	.ZN(n341));
   AOI22_X1 U356 (.A1(n346),
	.A2(n171),
	.B1(n291),
	.B2(n298),
	.ZN(n345));
   NOR2_X1 U357 (.A1(n45),
	.A2(n170),
	.ZN(n298));
   OAI221_X1 U358 (.A(n347),
	.B1(n305),
	.B2(n332),
	.C1(n304),
	.C2(n319),
	.ZN(n346));
   INV_X1 U359 (.A(n348),
	.ZN(n347));
   MUX2_X1 U360 (.A(n349),
	.B(n350),
	.S(ALU_OPB[2]),
	.Z(n348));
   NOR2_X1 U361 (.A1(n320),
	.A2(FE_DBTN13_ALU_OPA_28),
	.ZN(n350));
   OAI22_X1 U362 (.A1(n351),
	.A2(n352),
	.B1(n320),
	.B2(FE_DBTN11_ALU_OPA_24),
	.ZN(n349));
   MUX2_X1 U363 (.A(FE_DBTN12_ALU_OPA_26),
	.B(FE_DBTN14_ALU_OPA_30),
	.S(ALU_OPB[2]),
	.Z(n319));
   MUX2_X1 U364 (.A(n356),
	.B(n278),
	.S(ALU_OPB[2]),
	.Z(n332));
   NAND4_X1 U365 (.A1(n357),
	.A2(n358),
	.A3(n359),
	.A4(n360),
	.ZN(ALU_OUT[23]));
   OAI211_X1 U366 (.A(n171),
	.B(n307),
	.C1(n361),
	.C2(n362),
	.ZN(n360));
   INV_X1 U367 (.A(n344),
	.ZN(n307));
   OAI221_X1 U368 (.A(n366),
	.B1(FE_DBTN11_ALU_OPA_24),
	.B2(n363),
	.C1(n364),
	.C2(n365),
	.ZN(n362));
   AOI22_X1 U369 (.A1(n367),
	.A2(ALU_OPA[26]),
	.B1(n368),
	.B2(ALU_OPA[25]),
	.ZN(n366));
   OAI221_X1 U370 (.A(n371),
	.B1(FE_DBTN13_ALU_OPA_28),
	.B2(n369),
	.C1(n352),
	.C2(n370),
	.ZN(n361));
   AOI22_X1 U371 (.A1(n372),
	.A2(ALU_OPA[29]),
	.B1(n373),
	.B2(FE_OFN116_ALU_OPA_30),
	.ZN(n371));
   OAI21_X1 U372 (.A(n9),
	.B1(n374),
	.B2(n344),
	.ZN(n359));
   NAND2_X1 U373 (.A1(N695),
	.A2(FE_OFN34_n198),
	.ZN(n358));
   MUX2_X1 U374 (.A(n375),
	.B(n376),
	.S(ALU_OPB[23]),
	.Z(n357));
   MUX2_X1 U375 (.A(n4),
	.B(n201),
	.S(FE_OFN118_ALU_OPA_23),
	.Z(n376));
   NAND2_X1 U376 (.A1(FE_OFN118_ALU_OPA_23),
	.A2(FE_DBTN4_n4),
	.ZN(n375));
   NAND4_X1 U377 (.A1(n377),
	.A2(n378),
	.A3(n379),
	.A4(n380),
	.ZN(ALU_OUT[22]));
   OAI211_X1 U378 (.A(n171),
	.B(n383),
	.C1(n381),
	.C2(n382),
	.ZN(n380));
   INV_X1 U379 (.A(n384),
	.ZN(n383));
   OAI221_X1 U380 (.A(n386),
	.B1(n363),
	.B2(n365),
	.C1(n364),
	.C2(FE_DBTN10_ALU_OPA_22),
	.ZN(n382));
   AOI22_X1 U381 (.A1(n367),
	.A2(ALU_OPA[25]),
	.B1(n368),
	.B2(FE_OFN117_ALU_OPA_24),
	.ZN(n386));
   OAI221_X1 U382 (.A(n387),
	.B1(n352),
	.B2(n369),
	.C1(FE_DBTN12_ALU_OPA_26),
	.C2(n370),
	.ZN(n381));
   AOI222_X1 U383 (.A1(n373),
	.A2(ALU_OPA[29]),
	.B1(n374),
	.B2(FE_OFN116_ALU_OPA_30),
	.C1(n372),
	.C2(ALU_OPA[28]),
	.ZN(n387));
   OAI21_X1 U384 (.A(n9),
	.B1(n388),
	.B2(n384),
	.ZN(n379));
   OAI21_X1 U385 (.A(n390),
	.B1(FE_OFN115_ALU_OPB_0),
	.B2(n389),
	.ZN(n384));
   NAND2_X1 U386 (.A1(N694),
	.A2(FE_OFN34_n198),
	.ZN(n378));
   MUX2_X1 U387 (.A(n391),
	.B(n392),
	.S(ALU_OPB[22]),
	.Z(n377));
   MUX2_X1 U388 (.A(n4),
	.B(n201),
	.S(ALU_OPA[22]),
	.Z(n392));
   NAND2_X1 U389 (.A1(ALU_OPA[22]),
	.A2(FE_DBTN4_n4),
	.ZN(n391));
   NAND4_X1 U390 (.A1(n393),
	.A2(n394),
	.A3(n395),
	.A4(n396),
	.ZN(ALU_OUT[21]));
   OAI211_X1 U391 (.A(n390),
	.B(n171),
	.C1(n397),
	.C2(n398),
	.ZN(n396));
   OAI221_X1 U392 (.A(n401),
	.B1(FE_DBTN14_ALU_OPA_30),
	.B2(n399),
	.C1(n364),
	.C2(n400),
	.ZN(n398));
   AOI222_X1 U393 (.A1(ALU_OPA[22]),
	.A2(n402),
	.B1(n367),
	.B2(FE_OFN117_ALU_OPA_24),
	.C1(FE_OFN118_ALU_OPA_23),
	.C2(n368),
	.ZN(n401));
   OAI221_X1 U394 (.A(n403),
	.B1(FE_DBTN12_ALU_OPA_26),
	.B2(n369),
	.C1(n356),
	.C2(n370),
	.ZN(n397));
   AOI222_X1 U395 (.A1(n373),
	.A2(ALU_OPA[28]),
	.B1(n374),
	.B2(ALU_OPA[29]),
	.C1(n372),
	.C2(ALU_OPA[27]),
	.ZN(n403));
   INV_X1 U396 (.A(n404),
	.ZN(n395));
   AOI21_X1 U397 (.A(n170),
	.B1(n390),
	.B2(n405),
	.ZN(n404));
   OAI21_X1 U398 (.A(n344),
	.B1(n406),
	.B2(n284),
	.ZN(n390));
   NAND2_X1 U399 (.A1(n210),
	.A2(n389),
	.ZN(n344));
   NAND2_X1 U400 (.A1(N334),
	.A2(N331),
	.ZN(n284));
   INV_X1 U401 (.A(N332),
	.ZN(n406));
   NAND2_X1 U402 (.A1(N693),
	.A2(FE_OFN34_n198),
	.ZN(n394));
   MUX2_X1 U403 (.A(n407),
	.B(n408),
	.S(ALU_OPB[21]),
	.Z(n393));
   MUX2_X1 U404 (.A(n4),
	.B(n201),
	.S(ALU_OPA[21]),
	.Z(n408));
   NAND2_X1 U405 (.A1(ALU_OPA[21]),
	.A2(FE_DBTN4_n4),
	.ZN(n407));
   NAND4_X1 U406 (.A1(n409),
	.A2(n410),
	.A3(n411),
	.A4(n412),
	.ZN(ALU_OUT[20]));
   OAI211_X1 U407 (.A(n171),
	.B(n415),
	.C1(n413),
	.C2(n414),
	.ZN(n412));
   OAI221_X1 U408 (.A(n417),
	.B1(n364),
	.B2(FE_DBTN9_ALU_OPA_20),
	.C1(FE_DBTN14_ALU_OPA_30),
	.C2(n405),
	.ZN(n414));
   AOI222_X1 U409 (.A1(n388),
	.A2(ALU_OPA[29]),
	.B1(ALU_OPA[22]),
	.B2(n368),
	.C1(ALU_OPA[21]),
	.C2(n402),
	.ZN(n417));
   OAI211_X1 U410 (.A(n419),
	.B(n420),
	.C1(n418),
	.C2(n365),
	.ZN(n413));
   AOI222_X1 U411 (.A1(n373),
	.A2(ALU_OPA[27]),
	.B1(n374),
	.B2(ALU_OPA[28]),
	.C1(n372),
	.C2(ALU_OPA[26]),
	.ZN(n420));
   AOI22_X1 U412 (.A1(n421),
	.A2(ALU_OPA[25]),
	.B1(n422),
	.B2(FE_OFN117_ALU_OPA_24),
	.ZN(n419));
   INV_X1 U413 (.A(n423),
	.ZN(n411));
   AOI21_X1 U414 (.A(n170),
	.B1(n424),
	.B2(n415),
	.ZN(n423));
   INV_X1 U415 (.A(n425),
	.ZN(n415));
   OAI21_X1 U416 (.A(n426),
	.B1(n209),
	.B2(n389),
	.ZN(n425));
   NAND2_X1 U417 (.A1(N692),
	.A2(FE_OFN34_n198),
	.ZN(n410));
   MUX2_X1 U418 (.A(n427),
	.B(n428),
	.S(ALU_OPB[20]),
	.Z(n409));
   MUX2_X1 U419 (.A(n4),
	.B(n201),
	.S(ALU_OPA[20]),
	.Z(n428));
   NAND2_X1 U420 (.A1(ALU_OPA[20]),
	.A2(FE_DBTN4_n4),
	.ZN(n427));
   NAND3_X1 U421 (.A1(n429),
	.A2(n430),
	.A3(n431),
	.ZN(ALU_OUT[1]));
   MUX2_X1 U422 (.A(n170),
	.B(n432),
	.S(n433),
	.Z(n431));
   NAND2_X1 U423 (.A1(N665),
	.A2(n171),
	.ZN(n432));
   NAND2_X1 U424 (.A1(N673),
	.A2(FE_OFN34_n198),
	.ZN(n430));
   MUX2_X1 U425 (.A(n434),
	.B(n435),
	.S(ALU_OPB[1]),
	.Z(n429));
   MUX2_X1 U426 (.A(n4),
	.B(n201),
	.S(ALU_OPA[1]),
	.Z(n435));
   NAND2_X1 U427 (.A1(ALU_OPA[1]),
	.A2(FE_OFN42_FE_DBTN4_n4),
	.ZN(n434));
   NAND2_X1 U428 (.A1(n436),
	.A2(n437),
	.ZN(ALU_OUT[19]));
   MUX2_X1 U429 (.A(n438),
	.B(n439),
	.S(ALU_OPB[19]),
	.Z(n437));
   MUX2_X1 U430 (.A(n4),
	.B(n201),
	.S(ALU_OPA[19]),
	.Z(n439));
   NAND2_X1 U431 (.A1(ALU_OPA[19]),
	.A2(FE_OFN42_FE_DBTN4_n4),
	.ZN(n438));
   AOI21_X1 U432 (.A(n440),
	.B1(N691),
	.B2(FE_OFN34_n198),
	.ZN(n436));
   MUX2_X1 U433 (.A(n9),
	.B(n441),
	.S(n426),
	.Z(n440));
   NOR2_X1 U434 (.A1(n317),
	.A2(n442),
	.ZN(n426));
   OAI22_X1 U435 (.A1(n443),
	.A2(n10),
	.B1(n320),
	.B2(n444),
	.ZN(n441));
   NOR4_X1 U436 (.A1(n445),
	.A2(n446),
	.A3(n447),
	.A4(n448),
	.ZN(n443));
   OAI222_X1 U437 (.A1(n278),
	.A2(n405),
	.B1(n364),
	.B2(n142),
	.C1(FE_DBTN14_ALU_OPA_30),
	.C2(n424),
	.ZN(n448));
   OAI222_X1 U438 (.A1(n363),
	.A2(FE_DBTN9_ALU_OPA_20),
	.B1(n449),
	.B2(n400),
	.C1(FE_DBTN13_ALU_OPA_28),
	.C2(n399),
	.ZN(n447));
   OAI222_X1 U439 (.A1(n370),
	.A2(n365),
	.B1(FE_DBTN11_ALU_OPA_24),
	.B2(n369),
	.C1(n418),
	.C2(FE_DBTN10_ALU_OPA_22),
	.ZN(n446));
   OAI222_X1 U440 (.A1(n356),
	.A2(n450),
	.B1(n352),
	.B2(n451),
	.C1(FE_DBTN12_ALU_OPA_26),
	.C2(n452),
	.ZN(n445));
   NAND2_X1 U441 (.A1(n453),
	.A2(n454),
	.ZN(ALU_OUT[18]));
   MUX2_X1 U442 (.A(n455),
	.B(n456),
	.S(ALU_OPB[18]),
	.Z(n454));
   MUX2_X1 U443 (.A(n4),
	.B(n201),
	.S(FE_OFN119_ALU_OPA_18),
	.Z(n456));
   NAND2_X1 U444 (.A1(FE_OFN119_ALU_OPA_18),
	.A2(FE_OFN42_FE_DBTN4_n4),
	.ZN(n455));
   AOI21_X1 U445 (.A(n457),
	.B1(N690),
	.B2(FE_OFN34_n198),
	.ZN(n453));
   MUX2_X1 U446 (.A(n9),
	.B(n458),
	.S(n459),
	.Z(n457));
   AOI21_X1 U447 (.A(n460),
	.B1(n442),
	.B2(FE_DBTN5_ALU_OPB_0),
	.ZN(n459));
   INV_X1 U448 (.A(n461),
	.ZN(n460));
   OAI22_X1 U449 (.A1(n462),
	.A2(n10),
	.B1(n305),
	.B2(n444),
	.ZN(n458));
   NOR4_X1 U450 (.A1(n463),
	.A2(n464),
	.A3(n465),
	.A4(n466),
	.ZN(n462));
   OAI222_X1 U451 (.A1(FE_DBTN13_ALU_OPA_28),
	.A2(n405),
	.B1(n364),
	.B2(FE_DBTN8_ALU_OPA_18),
	.C1(n278),
	.C2(n424),
	.ZN(n466));
   OAI222_X1 U452 (.A1(n363),
	.A2(n142),
	.B1(n449),
	.B2(FE_DBTN9_ALU_OPA_20),
	.C1(n352),
	.C2(n399),
	.ZN(n465));
   OAI222_X1 U453 (.A1(n370),
	.A2(FE_DBTN10_ALU_OPA_22),
	.B1(n369),
	.B2(n365),
	.C1(n418),
	.C2(n400),
	.ZN(n464));
   OAI221_X1 U455 (.A(n470),
	.B1(n468),
	.B2(n469),
	.C1(FE_DBTN12_ALU_OPA_26),
	.C2(n451),
	.ZN(n463));
   AOI22_X1 U456 (.A1(n372),
	.A2(FE_OFN117_ALU_OPA_24),
	.B1(n373),
	.B2(ALU_OPA[25]),
	.ZN(n470));
   NAND2_X1 U457 (.A1(n299),
	.A2(FE_OFN116_ALU_OPA_30),
	.ZN(n469));
   NAND3_X1 U458 (.A1(n471),
	.A2(n472),
	.A3(n473),
	.ZN(ALU_OUT[17]));
   MUX2_X1 U459 (.A(n170),
	.B(n474),
	.S(n461),
	.Z(n473));
   AOI21_X1 U460 (.A(n317),
	.B1(n232),
	.B2(n442),
	.ZN(n461));
   NAND2_X1 U461 (.A1(n171),
	.A2(n475),
	.ZN(n474));
   NAND4_X1 U462 (.A1(n476),
	.A2(n477),
	.A3(n478),
	.A4(n479),
	.ZN(n475));
   AOI221_X1 U463 (.A(n482),
	.B1(n480),
	.B2(n481),
	.C1(n374),
	.C2(ALU_OPA[25]),
	.ZN(n479));
   OAI22_X1 U464 (.A1(FE_DBTN11_ALU_OPA_24),
	.A2(n452),
	.B1(n450),
	.B2(n365),
	.ZN(n482));
   INV_X1 U465 (.A(FE_OFN118_ALU_OPA_23),
	.ZN(n365));
   INV_X1 U466 (.A(n451),
	.ZN(n374));
   INV_X1 U467 (.A(n483),
	.ZN(n481));
   AOI21_X1 U468 (.A(n282),
	.B1(ALU_OPA[31]),
	.B2(n280),
	.ZN(n483));
   OAI22_X1 U469 (.A1(FE_DBTN14_ALU_OPA_30),
	.A2(n305),
	.B1(n320),
	.B2(n278),
	.ZN(n282));
   INV_X1 U470 (.A(ALU_OPA[29]),
	.ZN(n278));
   INV_X1 U471 (.A(n299),
	.ZN(n320));
   INV_X1 U472 (.A(n313),
	.ZN(n305));
   AOI222_X1 U474 (.A1(ALU_OPA[20]),
	.A2(n367),
	.B1(ALU_OPA[22]),
	.B2(n421),
	.C1(ALU_OPA[21]),
	.C2(n422),
	.ZN(n478));
   INV_X1 U475 (.A(n370),
	.ZN(n422));
   INV_X1 U476 (.A(n369),
	.ZN(n421));
   INV_X1 U477 (.A(n418),
	.ZN(n367));
   AOI222_X1 U478 (.A1(n388),
	.A2(ALU_OPA[26]),
	.B1(ALU_OPA[19]),
	.B2(n368),
	.C1(FE_OFN119_ALU_OPA_18),
	.C2(n402),
	.ZN(n477));
   INV_X1 U479 (.A(n363),
	.ZN(n402));
   INV_X1 U480 (.A(n449),
	.ZN(n368));
   INV_X1 U481 (.A(n399),
	.ZN(n388));
   INV_X1 U482 (.A(n484),
	.ZN(n476));
   OAI222_X1 U483 (.A1(n424),
	.A2(FE_DBTN13_ALU_OPA_28),
	.B1(n485),
	.B2(n364),
	.C1(n405),
	.C2(n352),
	.ZN(n484));
   NAND2_X1 U485 (.A1(N689),
	.A2(FE_OFN34_n198),
	.ZN(n472));
   MUX2_X1 U486 (.A(n486),
	.B(n487),
	.S(ALU_OPB[17]),
	.Z(n471));
   MUX2_X1 U487 (.A(n4),
	.B(n201),
	.S(ALU_OPA[17]),
	.Z(n487));
   NAND2_X1 U488 (.A1(ALU_OPA[17]),
	.A2(FE_OFN42_FE_DBTN4_n4),
	.ZN(n486));
   NAND2_X1 U489 (.A1(n488),
	.A2(n489),
	.ZN(ALU_OUT[16]));
   MUX2_X1 U490 (.A(n490),
	.B(n491),
	.S(ALU_OPB[16]),
	.Z(n489));
   MUX2_X1 U491 (.A(n4),
	.B(n201),
	.S(ALU_OPA[16]),
	.Z(n491));
   NAND2_X1 U492 (.A1(ALU_OPA[16]),
	.A2(FE_OFN42_FE_DBTN4_n4),
	.ZN(n490));
   AOI21_X1 U493 (.A(n492),
	.B1(N688),
	.B2(FE_OFN34_n198),
	.ZN(n488));
   MUX2_X1 U494 (.A(n9),
	.B(n493),
	.S(n494),
	.Z(n492));
   AOI21_X1 U495 (.A(n317),
	.B1(n442),
	.B2(n241),
	.ZN(n494));
   INV_X1 U496 (.A(n209),
	.ZN(n241));
   NAND2_X1 U497 (.A1(n232),
	.A2(FE_DBTN5_ALU_OPB_0),
	.ZN(n209));
   NOR2_X1 U498 (.A1(n389),
	.A2(N332),
	.ZN(n442));
   NAND2_X1 U499 (.A1(n329),
	.A2(n261),
	.ZN(n389));
   INV_X1 U500 (.A(N335),
	.ZN(n261));
   OAI22_X1 U501 (.A1(n495),
	.A2(n10),
	.B1(n351),
	.B2(n444),
	.ZN(n493));
   NAND2_X1 U502 (.A1(n480),
	.A2(n9),
	.ZN(n444));
   INV_X1 U503 (.A(n468),
	.ZN(n480));
   NOR4_X1 U504 (.A1(n496),
	.A2(n497),
	.A3(n498),
	.A4(n499),
	.ZN(n495));
   OAI222_X1 U505 (.A1(FE_DBTN12_ALU_OPA_26),
	.A2(n405),
	.B1(n364),
	.B2(FE_DBTN7_ALU_OPA_16),
	.C1(n352),
	.C2(n424),
	.ZN(n499));
   NAND2_X1 U506 (.A1(n501),
	.A2(n291),
	.ZN(n424));
   INV_X1 U507 (.A(ALU_OPA[27]),
	.ZN(n352));
   NAND2_X1 U509 (.A1(n502),
	.A2(n299),
	.ZN(n364));
   NAND2_X1 U510 (.A1(n501),
	.A2(n280),
	.ZN(n405));
   OAI222_X1 U512 (.A1(n363),
	.A2(n485),
	.B1(n449),
	.B2(FE_DBTN8_ALU_OPA_18),
	.C1(n356),
	.C2(n399),
	.ZN(n498));
   NAND2_X1 U513 (.A1(n501),
	.A2(n313),
	.ZN(n399));
   INV_X1 U514 (.A(ALU_OPA[25]),
	.ZN(n356));
   NAND2_X1 U516 (.A1(n502),
	.A2(n280),
	.ZN(n449));
   INV_X1 U517 (.A(ALU_OPA[17]),
	.ZN(n485));
   NAND2_X1 U518 (.A1(n502),
	.A2(n313),
	.ZN(n363));
   OAI222_X1 U519 (.A1(n370),
	.A2(FE_DBTN9_ALU_OPA_20),
	.B1(n369),
	.B2(n400),
	.C1(n418),
	.C2(n142),
	.ZN(n497));
   NAND2_X1 U520 (.A1(n502),
	.A2(n291),
	.ZN(n418));
   NOR2_X1 U521 (.A1(ALU_OPB[3]),
	.A2(ALU_OPB[2]),
	.ZN(n502));
   INV_X1 U522 (.A(ALU_OPA[21]),
	.ZN(n400));
   NAND2_X1 U523 (.A1(n503),
	.A2(n313),
	.ZN(n369));
   NAND2_X1 U525 (.A1(n503),
	.A2(n299),
	.ZN(n370));
   OAI221_X1 U526 (.A(n504),
	.B1(n289),
	.B2(n468),
	.C1(FE_DBTN11_ALU_OPA_24),
	.C2(n451),
	.ZN(n496));
   AOI22_X1 U527 (.A1(ALU_OPA[22]),
	.A2(n372),
	.B1(FE_OFN118_ALU_OPA_23),
	.B2(n373),
	.ZN(n504));
   INV_X1 U528 (.A(n452),
	.ZN(n373));
   NAND2_X1 U529 (.A1(n503),
	.A2(n291),
	.ZN(n452));
   INV_X1 U530 (.A(n351),
	.ZN(n291));
   NAND2_X1 U531 (.A1(ALU_OPB[1]),
	.A2(FE_OFN115_ALU_OPB_0),
	.ZN(n351));
   INV_X1 U532 (.A(n450),
	.ZN(n372));
   NAND2_X1 U533 (.A1(n503),
	.A2(n280),
	.ZN(n450));
   NOR2_X1 U534 (.A1(n45),
	.A2(ALU_OPB[3]),
	.ZN(n503));
   NAND2_X1 U535 (.A1(n501),
	.A2(n299),
	.ZN(n451));
   NOR2_X1 U536 (.A1(FE_DBTN6_ALU_OPB_3),
	.A2(ALU_OPB[2]),
	.ZN(n501));
   NAND2_X1 U538 (.A1(ALU_OPB[2]),
	.A2(ALU_OPB[3]),
	.ZN(n468));
   AOI222_X1 U539 (.A1(ALU_OPA[29]),
	.A2(n313),
	.B1(n299),
	.B2(ALU_OPA[28]),
	.C1(FE_OFN116_ALU_OPA_30),
	.C2(n280),
	.ZN(n289));
   NAND2_X1 U540 (.A1(ALU_OPB[1]),
	.A2(FE_DBTN5_ALU_OPB_0),
	.ZN(n304));
   NOR2_X1 U541 (.A1(FE_OFN115_ALU_OPB_0),
	.A2(ALU_OPB[1]),
	.ZN(n299));
   NOR2_X1 U542 (.A1(FE_DBTN5_ALU_OPB_0),
	.A2(ALU_OPB[1]),
	.ZN(n313));
   NAND3_X1 U543 (.A1(n505),
	.A2(n506),
	.A3(n507),
	.ZN(ALU_OUT[15]));
   MUX2_X1 U544 (.A(n508),
	.B(n170),
	.S(n317),
	.Z(n507));
   NAND2_X1 U545 (.A1(N591),
	.A2(n171),
	.ZN(n508));
   NAND2_X1 U546 (.A1(N687),
	.A2(FE_OFN34_n198),
	.ZN(n506));
   MUX2_X1 U547 (.A(n509),
	.B(n510),
	.S(ALU_OPB[15]),
	.Z(n505));
   MUX2_X1 U548 (.A(n4),
	.B(n201),
	.S(ALU_OPA[15]),
	.Z(n510));
   NAND2_X1 U549 (.A1(ALU_OPA[15]),
	.A2(FE_OFN42_FE_DBTN4_n4),
	.ZN(n509));
   NAND3_X1 U550 (.A1(n511),
	.A2(n512),
	.A3(n513),
	.ZN(ALU_OUT[14]));
   MUX2_X1 U551 (.A(n514),
	.B(n170),
	.S(n515),
	.Z(n513));
   AOI21_X1 U552 (.A(n210),
	.B1(n263),
	.B2(N332),
	.ZN(n515));
   INV_X1 U553 (.A(n317),
	.ZN(n210));
   NAND2_X1 U554 (.A1(N613),
	.A2(n171),
	.ZN(n514));
   NAND2_X1 U555 (.A1(N686),
	.A2(FE_OFN34_n198),
	.ZN(n512));
   MUX2_X1 U556 (.A(n516),
	.B(n517),
	.S(ALU_OPB[14]),
	.Z(n511));
   MUX2_X1 U557 (.A(n4),
	.B(n201),
	.S(FE_OFN120_ALU_OPA_14),
	.Z(n517));
   NAND2_X1 U558 (.A1(FE_OFN120_ALU_OPA_14),
	.A2(FE_OFN42_FE_DBTN4_n4),
	.ZN(n516));
   NAND3_X1 U559 (.A1(n518),
	.A2(n519),
	.A3(n520),
	.ZN(ALU_OUT[13]));
   MUX2_X1 U560 (.A(n170),
	.B(n521),
	.S(n522),
	.Z(n520));
   NAND2_X1 U561 (.A1(N617),
	.A2(n171),
	.ZN(n521));
   NAND2_X1 U562 (.A1(N685),
	.A2(FE_OFN34_n198),
	.ZN(n519));
   MUX2_X1 U563 (.A(n523),
	.B(n524),
	.S(ALU_OPB[13]),
	.Z(n518));
   MUX2_X1 U564 (.A(n4),
	.B(n201),
	.S(ALU_OPA[13]),
	.Z(n524));
   NAND2_X1 U565 (.A1(ALU_OPA[13]),
	.A2(FE_OFN42_FE_DBTN4_n4),
	.ZN(n523));
   NAND3_X1 U566 (.A1(n525),
	.A2(n526),
	.A3(n527),
	.ZN(ALU_OUT[12]));
   MUX2_X1 U567 (.A(n528),
	.B(n170),
	.S(n529),
	.Z(n527));
   AOI21_X1 U568 (.A(n522),
	.B1(n330),
	.B2(FE_OFN115_ALU_OPB_0),
	.ZN(n529));
   OAI21_X1 U569 (.A(n317),
	.B1(n232),
	.B2(n283),
	.ZN(n522));
   INV_X1 U570 (.A(n283),
	.ZN(n330));
   NAND2_X1 U571 (.A1(N621),
	.A2(n171),
	.ZN(n528));
   NAND2_X1 U572 (.A1(N684),
	.A2(FE_OFN34_n198),
	.ZN(n526));
   MUX2_X1 U573 (.A(n530),
	.B(n531),
	.S(ALU_OPB[12]),
	.Z(n525));
   MUX2_X1 U574 (.A(n4),
	.B(n201),
	.S(FE_OFN122_ALU_OPA_12),
	.Z(n531));
   NAND2_X1 U575 (.A1(FE_OFN122_ALU_OPA_12),
	.A2(FE_OFN42_FE_DBTN4_n4),
	.ZN(n530));
   NAND3_X1 U576 (.A1(n532),
	.A2(n533),
	.A3(n534),
	.ZN(ALU_OUT[11]));
   MUX2_X1 U577 (.A(n170),
	.B(n535),
	.S(n194),
	.Z(n534));
   NAND2_X1 U578 (.A1(N625),
	.A2(n171),
	.ZN(n535));
   NAND2_X1 U579 (.A1(N683),
	.A2(FE_OFN34_n198),
	.ZN(n533));
   MUX2_X1 U580 (.A(n536),
	.B(n537),
	.S(ALU_OPB[11]),
	.Z(n532));
   MUX2_X1 U581 (.A(n4),
	.B(n201),
	.S(ALU_OPA[11]),
	.Z(n537));
   NAND2_X1 U582 (.A1(ALU_OPA[11]),
	.A2(FE_OFN42_FE_DBTN4_n4),
	.ZN(n536));
   NAND3_X1 U583 (.A1(n538),
	.A2(n539),
	.A3(n540),
	.ZN(ALU_OUT[10]));
   MUX2_X1 U584 (.A(n541),
	.B(n170),
	.S(n542),
	.Z(n540));
   NOR2_X1 U585 (.A1(n263),
	.A2(n194),
	.ZN(n542));
   NAND2_X1 U586 (.A1(n317),
	.A2(n283),
	.ZN(n194));
   NAND2_X1 U587 (.A1(N333),
	.A2(N332),
	.ZN(n283));
   NOR3_X1 U588 (.A1(n232),
	.A2(n329),
	.A3(FE_DBTN5_ALU_OPB_0),
	.ZN(n263));
   NAND2_X1 U589 (.A1(N629),
	.A2(n171),
	.ZN(n541));
   NAND2_X1 U590 (.A1(N682),
	.A2(FE_OFN34_n198),
	.ZN(n539));
   MUX2_X1 U591 (.A(n543),
	.B(n544),
	.S(ALU_OPB[10]),
	.Z(n538));
   MUX2_X1 U592 (.A(n4),
	.B(n201),
	.S(FE_OFN121_ALU_OPA_10),
	.Z(n544));
   NAND2_X1 U593 (.A1(FE_OFN121_ALU_OPA_10),
	.A2(FE_OFN42_FE_DBTN4_n4),
	.ZN(n543));
   NAND4_X1 U594 (.A1(n545),
	.A2(n546),
	.A3(n547),
	.A4(n548),
	.ZN(ALU_OUT[0]));
   NAND4_X1 U595 (.A1(N671),
	.A2(OP[2]),
	.A3(n549),
	.A4(n550),
	.ZN(n548));
   NAND2_X1 U596 (.A1(N672),
	.A2(FE_OFN34_n198),
	.ZN(n547));
   XNOR2_X1 U597 (.A(n551),
	.B(OP[2]),
	.ZN(n198));
   NAND2_X1 U598 (.A1(n550),
	.A2(n549),
	.ZN(n551));
   MUX2_X1 U599 (.A(n552),
	.B(n553),
	.S(FE_OFN115_ALU_OPB_0),
	.Z(n546));
   MUX2_X1 U600 (.A(n4),
	.B(n201),
	.S(ALU_OPA[0]),
	.Z(n553));
   INV_X1 U601 (.A(n277),
	.ZN(n201));
   NOR3_X1 U602 (.A1(OP[1]),
	.A2(OP[2]),
	.A3(n549),
	.ZN(n277));
   NAND2_X1 U603 (.A1(ALU_OPA[0]),
	.A2(FE_OFN42_FE_DBTN4_n4),
	.ZN(n552));
   MUX2_X1 U604 (.A(n554),
	.B(n170),
	.S(n555),
	.Z(n545));
   NOR2_X1 U605 (.A1(FE_OFN115_ALU_OPB_0),
	.A2(n433),
	.ZN(n555));
   NAND2_X1 U606 (.A1(n233),
	.A2(n232),
	.ZN(n433));
   INV_X1 U607 (.A(N331),
	.ZN(n232));
   NOR2_X1 U608 (.A1(n224),
	.A2(N332),
	.ZN(n233));
   NAND2_X1 U609 (.A1(n317),
	.A2(n329),
	.ZN(n224));
   INV_X1 U610 (.A(N333),
	.ZN(n329));
   NAND2_X1 U611 (.A1(N669),
	.A2(n171),
	.ZN(n554));
   INV_X1 U612 (.A(OP[0]),
	.ZN(n549));
   INV_X1 U613 (.A(OP[1]),
	.ZN(n550));
endmodule

module exe_unit (
	clk, 
	rst, 
	en, 
	RF_OUT1, 
	RF_OUT2, 
	PC, 
	IMM, 
	EXE_MEM_IN, 
	MEM_WB_IN, 
	RD_IN, 
	RS1_IN, 
	RS2_IN, 
	ALU_OP, 
	ALU_OPA_SEL, 
	ALU_OPB_SEL, 
	ALU_OUT, 
	MEM_DATA, 
	RD_OUT, 
	RS1_OUT, 
	RS2_OUT);
   input clk;
   input rst;
   input en;
   input [31:0] RF_OUT1;
   input [31:0] RF_OUT2;
   input [31:0] PC;
   input [31:0] IMM;
   input [31:0] EXE_MEM_IN;
   input [31:0] MEM_WB_IN;
   input [4:0] RD_IN;
   input [4:0] RS1_IN;
   input [4:0] RS2_IN;
   input [2:0] ALU_OP;
   input [2:0] ALU_OPA_SEL;
   input [2:0] ALU_OPB_SEL;
   output [31:0] ALU_OUT;
   output [31:0] MEM_DATA;
   output [4:0] RD_OUT;
   output [4:0] RS1_OUT;
   output [4:0] RS2_OUT;

   // Internal wires
   wire FE_OFN104_n391;
   wire FE_OFN100_n391;
   wire FE_OFN95_n429;
   wire FE_OFN94_n430;
   wire FE_OFN91_n432;
   wire FE_OFN90_n432;
   wire FE_OFN45_n246;
   wire FE_OFN44_n246;
   wire FE_OFN43_n246;
   wire FE_OFN40_ALU_OPA_SEL_c_2;
   wire FE_OFN39_ALU_OPA_SEL_c_2;
   wire FE_OFN28_n394;
   wire FE_OFN27_n394;
   wire FE_OFN26_n394;
   wire FE_OFN25_n394;
   wire FE_OFN24_n394;
   wire FE_OFN23_n394;
   wire FE_OFN22_n393;
   wire FE_OFN20_n393;
   wire FE_OFN19_n393;
   wire FE_OFN2_n247;
   wire FE_OFN1_n247;
   wire FE_OFN0_n247;
   wire FE_DBTN3_ALU_OPA_SEL_c_2;
   wire FE_DBTN0_n37;
   wire n532;
   wire n12;
   wire n14;
   wire n16;
   wire n18;
   wire n20;
   wire n22;
   wire n24;
   wire n26;
   wire n28;
   wire n30;
   wire n32;
   wire n34;
   wire n36;
   wire n38;
   wire n40;
   wire n42;
   wire n44;
   wire n46;
   wire n48;
   wire n50;
   wire n52;
   wire n54;
   wire n56;
   wire n58;
   wire n60;
   wire n62;
   wire n64;
   wire n66;
   wire n68;
   wire n70;
   wire n72;
   wire n74;
   wire n245;
   wire n246;
   wire n247;
   wire n248;
   wire n249;
   wire n250;
   wire n251;
   wire n252;
   wire n253;
   wire n254;
   wire n255;
   wire n256;
   wire n257;
   wire n258;
   wire n259;
   wire n260;
   wire n261;
   wire n262;
   wire n263;
   wire n264;
   wire n265;
   wire n266;
   wire n267;
   wire n268;
   wire n269;
   wire n270;
   wire n271;
   wire n272;
   wire n273;
   wire n274;
   wire n275;
   wire n276;
   wire n277;
   wire n278;
   wire n279;
   wire n280;
   wire n281;
   wire n282;
   wire n283;
   wire n284;
   wire n285;
   wire n286;
   wire n287;
   wire n288;
   wire n289;
   wire n290;
   wire n291;
   wire n292;
   wire n293;
   wire n294;
   wire n295;
   wire n296;
   wire n297;
   wire n298;
   wire n299;
   wire n300;
   wire n301;
   wire n302;
   wire n303;
   wire n304;
   wire n305;
   wire n306;
   wire n307;
   wire n308;
   wire n309;
   wire n310;
   wire n311;
   wire n312;
   wire n313;
   wire n314;
   wire n315;
   wire n316;
   wire n317;
   wire n318;
   wire n319;
   wire n320;
   wire n321;
   wire n322;
   wire n323;
   wire n324;
   wire n325;
   wire n326;
   wire n327;
   wire n328;
   wire n329;
   wire n330;
   wire n331;
   wire n332;
   wire n333;
   wire n334;
   wire n335;
   wire n336;
   wire n337;
   wire n338;
   wire n339;
   wire n340;
   wire n341;
   wire n342;
   wire n343;
   wire n344;
   wire n345;
   wire n346;
   wire n347;
   wire n348;
   wire n349;
   wire n350;
   wire n351;
   wire n352;
   wire n353;
   wire n354;
   wire n355;
   wire n356;
   wire n357;
   wire n358;
   wire n359;
   wire n360;
   wire n361;
   wire n362;
   wire n363;
   wire n364;
   wire n365;
   wire n366;
   wire n367;
   wire n368;
   wire n369;
   wire n370;
   wire n371;
   wire n372;
   wire n373;
   wire n374;
   wire n375;
   wire n376;
   wire n377;
   wire n378;
   wire n379;
   wire n380;
   wire n381;
   wire n382;
   wire n383;
   wire n384;
   wire n385;
   wire n386;
   wire n387;
   wire n388;
   wire n389;
   wire n391;
   wire n392;
   wire n393;
   wire n394;
   wire n395;
   wire n396;
   wire n397;
   wire n398;
   wire n399;
   wire n400;
   wire n401;
   wire n402;
   wire n405;
   wire n406;
   wire n407;
   wire n408;
   wire n409;
   wire n410;
   wire n411;
   wire n412;
   wire n413;
   wire n414;
   wire n415;
   wire n416;
   wire n417;
   wire n418;
   wire n419;
   wire n420;
   wire n421;
   wire n422;
   wire n423;
   wire n424;
   wire n425;
   wire n426;
   wire n427;
   wire n428;
   wire n429;
   wire n430;
   wire n431;
   wire n432;
   wire n433;
   wire n434;
   wire n435;
   wire n436;
   wire n437;
   wire n438;
   wire n439;
   wire n440;
   wire n441;
   wire n442;
   wire n443;
   wire n444;
   wire n445;
   wire n446;
   wire n447;
   wire n448;
   wire n449;
   wire n450;
   wire n451;
   wire n452;
   wire n453;
   wire n454;
   wire n455;
   wire n456;
   wire n457;
   wire n458;
   wire n459;
   wire n460;
   wire n461;
   wire n462;
   wire n463;
   wire n1;
   wire n2;
   wire n3;
   wire n5;
   wire n6;
   wire n8;
   wire n9;
   wire n33;
   wire n55;
   wire n107;
   wire n108;
   wire n109;
   wire n110;
   wire n111;
   wire n112;
   wire n113;
   wire n114;
   wire n115;
   wire n116;
   wire n117;
   wire n118;
   wire n119;
   wire n120;
   wire n121;
   wire n122;
   wire n123;
   wire n124;
   wire n125;
   wire n126;
   wire n127;
   wire n128;
   wire n129;
   wire n130;
   wire n131;
   wire n132;
   wire n133;
   wire n134;
   wire n135;
   wire n136;
   wire n137;
   wire n138;
   wire n139;
   wire n140;
   wire n141;
   wire n142;
   wire n143;
   wire n144;
   wire n145;
   wire n146;
   wire n147;
   wire n148;
   wire n149;
   wire n150;
   wire n151;
   wire n152;
   wire n153;
   wire n154;
   wire n155;
   wire n156;
   wire n157;
   wire n158;
   wire n159;
   wire n160;
   wire n161;
   wire n162;
   wire n163;
   wire n164;
   wire n165;
   wire n166;
   wire n167;
   wire n168;
   wire n169;
   wire n170;
   wire n171;
   wire n172;
   wire n173;
   wire n174;
   wire n175;
   wire n176;
   wire n177;
   wire n178;
   wire n179;
   wire n180;
   wire n181;
   wire n182;
   wire n183;
   wire n184;
   wire n185;
   wire n186;
   wire n187;
   wire n188;
   wire n189;
   wire n190;
   wire n191;
   wire n192;
   wire n193;
   wire n194;
   wire n195;
   wire n196;
   wire n197;
   wire n198;
   wire n199;
   wire n200;
   wire n201;
   wire n202;
   wire n203;
   wire n204;
   wire n205;
   wire n206;
   wire n207;
   wire n208;
   wire n209;
   wire n210;
   wire n211;
   wire n212;
   wire n213;
   wire n214;
   wire n215;
   wire n216;
   wire n217;
   wire n218;
   wire n219;
   wire n220;
   wire n221;
   wire n222;
   wire n223;
   wire n224;
   wire n225;
   wire n226;
   wire n227;
   wire n228;
   wire n229;
   wire n230;
   wire n231;
   wire n232;
   wire n233;
   wire n234;
   wire n235;
   wire n236;
   wire n237;
   wire n238;
   wire n239;
   wire n240;
   wire n241;
   wire n242;
   wire n243;
   wire n244;
   wire n390;
   wire n403;
   wire n404;
   wire n464;
   wire n465;
   wire n466;
   wire n467;
   wire n468;
   wire n469;
   wire n470;
   wire n471;
   wire n472;
   wire n473;
   wire n474;
   wire n475;
   wire n476;
   wire n477;
   wire n478;
   wire n479;
   wire n480;
   wire n481;
   wire n482;
   wire n483;
   wire n484;
   wire n485;
   wire n486;
   wire n487;
   wire n488;
   wire n489;
   wire n490;
   wire n491;
   wire n492;
   wire n493;
   wire n494;
   wire n495;
   wire n496;
   wire n497;
   wire n498;
   wire n499;
   wire n500;
   wire n501;
   wire n502;
   wire n503;
   wire n504;
   wire n505;
   wire n506;
   wire n507;
   wire n508;
   wire n509;
   wire n510;
   wire n511;
   wire n512;
   wire n513;
   wire n514;
   wire n515;
   wire n516;
   wire n517;
   wire n518;
   wire n519;
   wire n520;
   wire n521;
   wire n522;
   wire n523;
   wire n524;
   wire n525;
   wire n526;
   wire n527;
   wire n528;
   wire n529;
   wire n530;
   wire n531;
   wire [31:0] ALU_OPA;
   wire [31:0] ALU_OPB;
   wire [31:0] currRF1;
   wire [31:0] currPC;
   wire [31:0] currIMM;

   BUF_X1 FE_OFC104_n391 (.A(FE_OFN100_n391),
	.Z(FE_OFN104_n391));
   BUF_X1 FE_OFC100_n391 (.A(n391),
	.Z(FE_OFN100_n391));
   BUF_X1 FE_OFC95_n429 (.A(n429),
	.Z(FE_OFN95_n429));
   BUF_X1 FE_OFC94_n430 (.A(n430),
	.Z(FE_OFN94_n430));
   BUF_X1 FE_OFC91_n432 (.A(FE_OFN90_n432),
	.Z(FE_OFN91_n432));
   BUF_X1 FE_OFC90_n432 (.A(n432),
	.Z(FE_OFN90_n432));
   CLKBUF_X3 FE_OFC45_n246 (.A(FE_OFN44_n246),
	.Z(FE_OFN45_n246));
   BUF_X1 FE_OFC44_n246 (.A(FE_OFN43_n246),
	.Z(FE_OFN44_n246));
   CLKBUF_X3 FE_OFC43_n246 (.A(n246),
	.Z(FE_OFN43_n246));
   BUF_X1 FE_OFC40_ALU_OPA_SEL_c_2 (.A(FE_OFN39_ALU_OPA_SEL_c_2),
	.Z(FE_OFN40_ALU_OPA_SEL_c_2));
   BUF_X1 FE_OFC39_ALU_OPA_SEL_c_2 (.A(ALU_OPA_SEL[2]),
	.Z(FE_OFN39_ALU_OPA_SEL_c_2));
   BUF_X1 FE_OFC28_n394 (.A(FE_OFN23_n394),
	.Z(FE_OFN28_n394));
   BUF_X1 FE_OFC27_n394 (.A(FE_OFN23_n394),
	.Z(FE_OFN27_n394));
   BUF_X1 FE_OFC26_n394 (.A(FE_OFN23_n394),
	.Z(FE_OFN26_n394));
   BUF_X1 FE_OFC25_n394 (.A(FE_OFN23_n394),
	.Z(FE_OFN25_n394));
   BUF_X1 FE_OFC24_n394 (.A(FE_OFN23_n394),
	.Z(FE_OFN24_n394));
   BUF_X1 FE_OFC23_n394 (.A(n394),
	.Z(FE_OFN23_n394));
   BUF_X1 FE_OFC22_n393 (.A(FE_OFN20_n393),
	.Z(FE_OFN22_n393));
   BUF_X1 FE_OFC20_n393 (.A(FE_OFN19_n393),
	.Z(FE_OFN20_n393));
   BUF_X1 FE_OFC19_n393 (.A(n393),
	.Z(FE_OFN19_n393));
   CLKBUF_X3 FE_OFC2_n247 (.A(FE_OFN1_n247),
	.Z(FE_OFN2_n247));
   BUF_X1 FE_OFC1_n247 (.A(FE_OFN0_n247),
	.Z(FE_OFN1_n247));
   CLKBUF_X3 FE_OFC0_n247 (.A(n247),
	.Z(FE_OFN0_n247));
   INV_X1 FE_DBTC3_ALU_OPA_SEL_c_2 (.A(ALU_OPA_SEL[2]),
	.ZN(FE_DBTN3_ALU_OPA_SEL_c_2));
   INV_X2 FE_DBTC0_n37 (.A(n8),
	.ZN(FE_DBTN0_n37));
   DFF_X1 currRS2_reg_4_ (.D(n237),
	.CK(clk),
	.Q(RS2_OUT[4]));
   DFF_X1 currRS2_reg_3_ (.D(n238),
	.CK(clk),
	.Q(RS2_OUT[3]));
   DFF_X1 currRS2_reg_2_ (.D(n239),
	.CK(clk),
	.Q(n532),
	.QN(n9));
   DFF_X1 currRS2_reg_1_ (.D(n240),
	.CK(clk),
	.Q(RS2_OUT[1]));
   DFF_X1 currRD_reg_4_ (.D(n242),
	.CK(clk),
	.Q(RD_OUT[4]));
   DFF_X1 currRD_reg_3_ (.D(n243),
	.CK(clk),
	.Q(RD_OUT[3]));
   DFF_X1 currRD_reg_2_ (.D(n244),
	.CK(clk),
	.Q(RD_OUT[2]));
   DFF_X1 currRD_reg_1_ (.D(n390),
	.CK(clk),
	.Q(RD_OUT[1]));
   DFF_X1 currRD_reg_0_ (.D(n403),
	.CK(clk),
	.Q(RD_OUT[0]));
   DFF_X1 currRF1_reg_31_ (.D(n107),
	.CK(clk),
	.Q(currRF1[31]),
	.QN(n12));
   DFF_X1 currRF1_reg_30_ (.D(n109),
	.CK(clk),
	.Q(currRF1[30]),
	.QN(n14));
   DFF_X1 currRF1_reg_29_ (.D(n111),
	.CK(clk),
	.Q(currRF1[29]),
	.QN(n16));
   DFF_X1 currRF1_reg_28_ (.D(n113),
	.CK(clk),
	.Q(currRF1[28]),
	.QN(n18));
   DFF_X1 currRF1_reg_27_ (.D(n115),
	.CK(clk),
	.Q(currRF1[27]),
	.QN(n20));
   DFF_X1 currRF1_reg_26_ (.D(n117),
	.CK(clk),
	.Q(currRF1[26]),
	.QN(n22));
   DFF_X1 currRF1_reg_25_ (.D(n119),
	.CK(clk),
	.Q(currRF1[25]),
	.QN(n24));
   DFF_X1 currRF1_reg_24_ (.D(n121),
	.CK(clk),
	.Q(currRF1[24]),
	.QN(n26));
   DFF_X1 currRF1_reg_23_ (.D(n123),
	.CK(clk),
	.Q(currRF1[23]),
	.QN(n28));
   DFF_X1 currRF1_reg_22_ (.D(n125),
	.CK(clk),
	.Q(currRF1[22]),
	.QN(n30));
   DFF_X1 currRF1_reg_21_ (.D(n127),
	.CK(clk),
	.Q(currRF1[21]),
	.QN(n32));
   DFF_X1 currRF1_reg_20_ (.D(n129),
	.CK(clk),
	.Q(currRF1[20]),
	.QN(n34));
   DFF_X1 currRF1_reg_19_ (.D(n131),
	.CK(clk),
	.Q(currRF1[19]),
	.QN(n36));
   DFF_X1 currRF1_reg_18_ (.D(n133),
	.CK(clk),
	.Q(currRF1[18]),
	.QN(n38));
   DFF_X1 currRF1_reg_17_ (.D(n135),
	.CK(clk),
	.Q(currRF1[17]),
	.QN(n40));
   DFF_X1 currRF1_reg_16_ (.D(n137),
	.CK(clk),
	.Q(currRF1[16]),
	.QN(n42));
   DFF_X1 currRF1_reg_15_ (.D(n139),
	.CK(clk),
	.Q(currRF1[15]),
	.QN(n44));
   DFF_X1 currRF1_reg_14_ (.D(n141),
	.CK(clk),
	.Q(currRF1[14]),
	.QN(n46));
   DFF_X1 currRF1_reg_13_ (.D(n143),
	.CK(clk),
	.Q(currRF1[13]),
	.QN(n48));
   DFF_X1 currRF1_reg_12_ (.D(n145),
	.CK(clk),
	.Q(currRF1[12]),
	.QN(n50));
   DFF_X1 currRF1_reg_11_ (.D(n147),
	.CK(clk),
	.Q(currRF1[11]),
	.QN(n52));
   DFF_X1 currRF1_reg_10_ (.D(n149),
	.CK(clk),
	.Q(currRF1[10]),
	.QN(n54));
   DFF_X1 currRF1_reg_9_ (.D(n151),
	.CK(clk),
	.Q(currRF1[9]),
	.QN(n56));
   DFF_X1 currRF1_reg_8_ (.D(n153),
	.CK(clk),
	.Q(currRF1[8]),
	.QN(n58));
   DFF_X1 currRF1_reg_7_ (.D(n155),
	.CK(clk),
	.Q(currRF1[7]),
	.QN(n60));
   DFF_X1 currRF1_reg_6_ (.D(n157),
	.CK(clk),
	.Q(currRF1[6]),
	.QN(n62));
   DFF_X1 currRF1_reg_5_ (.D(n159),
	.CK(clk),
	.Q(currRF1[5]),
	.QN(n64));
   DFF_X1 currRF1_reg_4_ (.D(n161),
	.CK(clk),
	.Q(currRF1[4]),
	.QN(n66));
   DFF_X1 currRF1_reg_3_ (.D(n163),
	.CK(clk),
	.Q(currRF1[3]),
	.QN(n68));
   DFF_X1 currRF1_reg_2_ (.D(n165),
	.CK(clk),
	.Q(currRF1[2]),
	.QN(n70));
   DFF_X1 currRF1_reg_1_ (.D(n167),
	.CK(clk),
	.Q(currRF1[1]),
	.QN(n72));
   DFF_X1 currRF1_reg_0_ (.D(n169),
	.CK(clk),
	.Q(currRF1[0]),
	.QN(n74));
   DFF_X1 currRF2_reg_31_ (.D(n108),
	.CK(clk),
	.Q(MEM_DATA[31]));
   DFF_X1 currRF2_reg_30_ (.D(n110),
	.CK(clk),
	.Q(MEM_DATA[30]));
   DFF_X1 currRF2_reg_29_ (.D(n112),
	.CK(clk),
	.Q(MEM_DATA[29]));
   DFF_X1 currRF2_reg_28_ (.D(n114),
	.CK(clk),
	.Q(MEM_DATA[28]));
   DFF_X1 currRF2_reg_27_ (.D(n116),
	.CK(clk),
	.Q(MEM_DATA[27]));
   DFF_X1 currRF2_reg_26_ (.D(n118),
	.CK(clk),
	.Q(MEM_DATA[26]));
   DFF_X1 currRF2_reg_25_ (.D(n120),
	.CK(clk),
	.Q(MEM_DATA[25]));
   DFF_X1 currRF2_reg_24_ (.D(n122),
	.CK(clk),
	.Q(MEM_DATA[24]));
   DFF_X1 currRF2_reg_23_ (.D(n124),
	.CK(clk),
	.Q(MEM_DATA[23]));
   DFF_X1 currRF2_reg_22_ (.D(n126),
	.CK(clk),
	.Q(MEM_DATA[22]));
   DFF_X1 currRF2_reg_21_ (.D(n128),
	.CK(clk),
	.Q(MEM_DATA[21]));
   DFF_X1 currRF2_reg_20_ (.D(n130),
	.CK(clk),
	.Q(MEM_DATA[20]));
   DFF_X1 currRF2_reg_19_ (.D(n132),
	.CK(clk),
	.Q(MEM_DATA[19]));
   DFF_X1 currRF2_reg_18_ (.D(n134),
	.CK(clk),
	.Q(MEM_DATA[18]));
   DFF_X1 currRF2_reg_17_ (.D(n136),
	.CK(clk),
	.Q(MEM_DATA[17]));
   DFF_X1 currRF2_reg_16_ (.D(n138),
	.CK(clk),
	.Q(MEM_DATA[16]));
   DFF_X1 currRF2_reg_15_ (.D(n140),
	.CK(clk),
	.Q(MEM_DATA[15]));
   DFF_X1 currRF2_reg_14_ (.D(n142),
	.CK(clk),
	.Q(MEM_DATA[14]));
   DFF_X1 currRF2_reg_13_ (.D(n144),
	.CK(clk),
	.Q(MEM_DATA[13]));
   DFF_X1 currRF2_reg_12_ (.D(n146),
	.CK(clk),
	.Q(MEM_DATA[12]));
   DFF_X1 currRF2_reg_11_ (.D(n148),
	.CK(clk),
	.Q(MEM_DATA[11]));
   DFF_X1 currRF2_reg_10_ (.D(n150),
	.CK(clk),
	.Q(MEM_DATA[10]));
   DFF_X1 currRF2_reg_9_ (.D(n152),
	.CK(clk),
	.Q(MEM_DATA[9]));
   DFF_X1 currRF2_reg_8_ (.D(n154),
	.CK(clk),
	.Q(MEM_DATA[8]));
   DFF_X1 currRF2_reg_7_ (.D(n156),
	.CK(clk),
	.Q(MEM_DATA[7]));
   DFF_X1 currRF2_reg_6_ (.D(n158),
	.CK(clk),
	.Q(MEM_DATA[6]));
   DFF_X1 currRF2_reg_5_ (.D(n160),
	.CK(clk),
	.Q(MEM_DATA[5]));
   DFF_X1 currRF2_reg_4_ (.D(n162),
	.CK(clk),
	.Q(MEM_DATA[4]));
   DFF_X1 currRF2_reg_3_ (.D(n164),
	.CK(clk),
	.Q(MEM_DATA[3]));
   DFF_X1 currRF2_reg_2_ (.D(n166),
	.CK(clk),
	.Q(MEM_DATA[2]));
   DFF_X1 currRF2_reg_1_ (.D(n168),
	.CK(clk),
	.Q(MEM_DATA[1]));
   DFF_X1 currRF2_reg_0_ (.D(n170),
	.CK(clk),
	.Q(MEM_DATA[0]));
   DFF_X1 currPC_reg_31_ (.D(n404),
	.CK(clk),
	.Q(currPC[31]));
   DFF_X1 currPC_reg_30_ (.D(n464),
	.CK(clk),
	.Q(currPC[30]));
   DFF_X1 currPC_reg_29_ (.D(n465),
	.CK(clk),
	.Q(currPC[29]));
   DFF_X1 currPC_reg_28_ (.D(n466),
	.CK(clk),
	.Q(currPC[28]));
   DFF_X1 currPC_reg_27_ (.D(n467),
	.CK(clk),
	.Q(currPC[27]));
   DFF_X1 currPC_reg_26_ (.D(n468),
	.CK(clk),
	.Q(currPC[26]));
   DFF_X1 currPC_reg_25_ (.D(n469),
	.CK(clk),
	.Q(currPC[25]));
   DFF_X1 currPC_reg_24_ (.D(n470),
	.CK(clk),
	.Q(currPC[24]));
   DFF_X1 currPC_reg_23_ (.D(n471),
	.CK(clk),
	.Q(currPC[23]));
   DFF_X1 currPC_reg_22_ (.D(n472),
	.CK(clk),
	.Q(currPC[22]));
   DFF_X1 currPC_reg_21_ (.D(n473),
	.CK(clk),
	.Q(currPC[21]));
   DFF_X1 currPC_reg_20_ (.D(n474),
	.CK(clk),
	.Q(currPC[20]));
   DFF_X1 currPC_reg_19_ (.D(n475),
	.CK(clk),
	.Q(currPC[19]));
   DFF_X1 currPC_reg_18_ (.D(n476),
	.CK(clk),
	.Q(currPC[18]));
   DFF_X1 currPC_reg_17_ (.D(n477),
	.CK(clk),
	.Q(currPC[17]));
   DFF_X1 currPC_reg_16_ (.D(n478),
	.CK(clk),
	.Q(currPC[16]));
   DFF_X1 currPC_reg_15_ (.D(n479),
	.CK(clk),
	.Q(currPC[15]));
   DFF_X1 currPC_reg_14_ (.D(n480),
	.CK(clk),
	.Q(currPC[14]));
   DFF_X1 currPC_reg_13_ (.D(n481),
	.CK(clk),
	.Q(currPC[13]));
   DFF_X1 currPC_reg_12_ (.D(n482),
	.CK(clk),
	.Q(currPC[12]));
   DFF_X1 currPC_reg_11_ (.D(n483),
	.CK(clk),
	.Q(currPC[11]));
   DFF_X1 currPC_reg_10_ (.D(n484),
	.CK(clk),
	.Q(currPC[10]));
   DFF_X1 currPC_reg_9_ (.D(n485),
	.CK(clk),
	.Q(currPC[9]));
   DFF_X1 currPC_reg_8_ (.D(n486),
	.CK(clk),
	.Q(currPC[8]));
   DFF_X1 currPC_reg_7_ (.D(n487),
	.CK(clk),
	.Q(currPC[7]));
   DFF_X1 currPC_reg_6_ (.D(n488),
	.CK(clk),
	.Q(currPC[6]));
   DFF_X1 currPC_reg_5_ (.D(n489),
	.CK(clk),
	.Q(currPC[5]));
   DFF_X1 currPC_reg_4_ (.D(n490),
	.CK(clk),
	.Q(currPC[4]));
   DFF_X1 currPC_reg_3_ (.D(n491),
	.CK(clk),
	.Q(currPC[3]));
   DFF_X1 currPC_reg_2_ (.D(n492),
	.CK(clk),
	.Q(currPC[2]));
   DFF_X1 currPC_reg_1_ (.D(n493),
	.CK(clk),
	.Q(currPC[1]));
   DFF_X1 currPC_reg_0_ (.D(n494),
	.CK(clk),
	.Q(currPC[0]));
   DFF_X1 currIMM_reg_31_ (.D(n495),
	.CK(clk),
	.Q(currIMM[31]));
   DFF_X1 currIMM_reg_30_ (.D(n496),
	.CK(clk),
	.Q(currIMM[30]));
   DFF_X1 currIMM_reg_29_ (.D(n497),
	.CK(clk),
	.Q(currIMM[29]));
   DFF_X1 currIMM_reg_28_ (.D(n498),
	.CK(clk),
	.Q(currIMM[28]));
   DFF_X1 currIMM_reg_27_ (.D(n499),
	.CK(clk),
	.Q(currIMM[27]));
   DFF_X1 currIMM_reg_26_ (.D(n500),
	.CK(clk),
	.Q(currIMM[26]));
   DFF_X1 currIMM_reg_25_ (.D(n501),
	.CK(clk),
	.Q(currIMM[25]));
   DFF_X1 currIMM_reg_24_ (.D(n502),
	.CK(clk),
	.Q(currIMM[24]));
   DFF_X1 currIMM_reg_23_ (.D(n503),
	.CK(clk),
	.Q(currIMM[23]));
   DFF_X1 currIMM_reg_22_ (.D(n504),
	.CK(clk),
	.Q(currIMM[22]));
   DFF_X1 currIMM_reg_21_ (.D(n505),
	.CK(clk),
	.Q(currIMM[21]));
   DFF_X1 currIMM_reg_20_ (.D(n506),
	.CK(clk),
	.Q(currIMM[20]));
   DFF_X1 currIMM_reg_19_ (.D(n507),
	.CK(clk),
	.Q(currIMM[19]));
   DFF_X1 currIMM_reg_18_ (.D(n508),
	.CK(clk),
	.Q(currIMM[18]));
   DFF_X1 currIMM_reg_17_ (.D(n509),
	.CK(clk),
	.Q(currIMM[17]));
   DFF_X1 currIMM_reg_16_ (.D(n510),
	.CK(clk),
	.Q(currIMM[16]));
   DFF_X1 currIMM_reg_15_ (.D(n511),
	.CK(clk),
	.Q(currIMM[15]));
   DFF_X1 currIMM_reg_14_ (.D(n512),
	.CK(clk),
	.Q(currIMM[14]));
   DFF_X1 currIMM_reg_13_ (.D(n513),
	.CK(clk),
	.Q(currIMM[13]));
   DFF_X1 currIMM_reg_12_ (.D(n514),
	.CK(clk),
	.Q(currIMM[12]));
   DFF_X1 currIMM_reg_11_ (.D(n515),
	.CK(clk),
	.Q(currIMM[11]));
   DFF_X1 currIMM_reg_10_ (.D(n516),
	.CK(clk),
	.Q(currIMM[10]));
   DFF_X1 currIMM_reg_9_ (.D(n517),
	.CK(clk),
	.Q(currIMM[9]));
   DFF_X1 currIMM_reg_8_ (.D(n518),
	.CK(clk),
	.Q(currIMM[8]));
   DFF_X1 currIMM_reg_7_ (.D(n519),
	.CK(clk),
	.Q(currIMM[7]));
   DFF_X1 currIMM_reg_6_ (.D(n520),
	.CK(clk),
	.Q(currIMM[6]));
   DFF_X1 currIMM_reg_5_ (.D(n521),
	.CK(clk),
	.Q(currIMM[5]));
   DFF_X1 currIMM_reg_4_ (.D(n522),
	.CK(clk),
	.Q(currIMM[4]));
   DFF_X1 currIMM_reg_3_ (.D(n523),
	.CK(clk),
	.Q(currIMM[3]));
   DFF_X1 currIMM_reg_2_ (.D(n524),
	.CK(clk),
	.Q(currIMM[2]));
   DFF_X1 currIMM_reg_1_ (.D(n525),
	.CK(clk),
	.Q(currIMM[1]));
   DFF_X1 currIMM_reg_0_ (.D(n526),
	.CK(clk),
	.Q(currIMM[0]));
   DFF_X1 currRS1_reg_4_ (.D(n527),
	.CK(clk),
	.Q(RS1_OUT[4]));
   DFF_X1 currRS1_reg_3_ (.D(n528),
	.CK(clk),
	.Q(RS1_OUT[3]));
   DFF_X1 currRS1_reg_1_ (.D(n530),
	.CK(clk),
	.Q(RS1_OUT[1]));
   NAND3_X1 U495 (.A1(FE_DBTN3_ALU_OPA_SEL_c_2),
	.A2(ALU_OPA_SEL[0]),
	.A3(ALU_OPA_SEL[1]),
	.ZN(n430));
   NAND3_X1 U496 (.A1(n171),
	.A2(FE_DBTN3_ALU_OPA_SEL_c_2),
	.A3(ALU_OPA_SEL[0]),
	.ZN(n429));
   alu_N32 alu_i (.OP(ALU_OP),
	.ALU_OPA(ALU_OPA),
	.ALU_OPB({ ALU_OPB[31],
		ALU_OPB[30],
		ALU_OPB[29],
		ALU_OPB[28],
		ALU_OPB[27],
		ALU_OPB[26],
		ALU_OPB[25],
		ALU_OPB[24],
		ALU_OPB[23],
		ALU_OPB[22],
		ALU_OPB[21],
		ALU_OPB[20],
		ALU_OPB[19],
		ALU_OPB[18],
		ALU_OPB[17],
		ALU_OPB[16],
		ALU_OPB[15],
		ALU_OPB[14],
		ALU_OPB[13],
		ALU_OPB[12],
		ALU_OPB[11],
		ALU_OPB[10],
		ALU_OPB[9],
		ALU_OPB[8],
		ALU_OPB[7],
		ALU_OPB[6],
		ALU_OPB[5],
		ALU_OPB[4],
		ALU_OPB[3],
		n33,
		ALU_OPB[1],
		ALU_OPB[0] }),
	.ALU_OUT(ALU_OUT));
   DFF_X1 currRS2_reg_0_ (.D(n241),
	.CK(clk),
	.Q(RS2_OUT[0]));
   DFF_X1 currRS1_reg_0_ (.D(n531),
	.CK(clk),
	.Q(RS1_OUT[0]));
   DFF_X1 currRS1_reg_2_ (.D(n529),
	.CK(clk),
	.Q(RS1_OUT[2]));
   OAI221_X4 U3 (.A(n443),
	.B1(n18),
	.B2(FE_OFN95_n429),
	.C1(n208),
	.C2(FE_OFN94_n430),
	.ZN(ALU_OPA[28]));
   OAI221_X4 U4 (.A(n442),
	.B1(n16),
	.B2(FE_OFN95_n429),
	.C1(n207),
	.C2(FE_OFN94_n430),
	.ZN(ALU_OPA[29]));
   OAI221_X2 U5 (.A(n439),
	.B1(n12),
	.B2(FE_OFN95_n429),
	.C1(n205),
	.C2(FE_OFN94_n430),
	.ZN(ALU_OPA[31]));
   OAI221_X4 U6 (.A(n444),
	.B1(n20),
	.B2(FE_OFN95_n429),
	.C1(n209),
	.C2(FE_OFN94_n430),
	.ZN(ALU_OPA[27]));
   OAI221_X2 U7 (.A(n445),
	.B1(n22),
	.B2(FE_OFN95_n429),
	.C1(n210),
	.C2(FE_OFN94_n430),
	.ZN(ALU_OPA[26]));
   OAI221_X4 U8 (.A(n446),
	.B1(n24),
	.B2(FE_OFN95_n429),
	.C1(n211),
	.C2(FE_OFN94_n430),
	.ZN(ALU_OPA[25]));
   OAI221_X4 U9 (.A(n449),
	.B1(n30),
	.B2(FE_OFN95_n429),
	.C1(n214),
	.C2(FE_OFN94_n430),
	.ZN(ALU_OPA[22]));
   OAI221_X2 U10 (.A(n451),
	.B1(n34),
	.B2(FE_OFN95_n429),
	.C1(n216),
	.C2(FE_OFN94_n430),
	.ZN(ALU_OPA[20]));
   OAI221_X2 U11 (.A(n453),
	.B1(n36),
	.B2(FE_OFN95_n429),
	.C1(n217),
	.C2(FE_OFN94_n430),
	.ZN(ALU_OPA[19]));
   OAI221_X4 U12 (.A(n455),
	.B1(n40),
	.B2(n429),
	.C1(n219),
	.C2(n430),
	.ZN(ALU_OPA[17]));
   OAI221_X4 U13 (.A(n456),
	.B1(n42),
	.B2(n429),
	.C1(n220),
	.C2(n430),
	.ZN(ALU_OPA[16]));
   OAI221_X4 U14 (.A(n457),
	.B1(n44),
	.B2(n429),
	.C1(n221),
	.C2(n430),
	.ZN(ALU_OPA[15]));
   OAI221_X4 U15 (.A(n459),
	.B1(n48),
	.B2(n429),
	.C1(n223),
	.C2(n430),
	.ZN(ALU_OPA[13]));
   OAI221_X4 U16 (.A(n461),
	.B1(n52),
	.B2(n429),
	.C1(n225),
	.C2(n430),
	.ZN(ALU_OPA[11]));
   OAI221_X4 U18 (.A(n450),
	.B1(n32),
	.B2(FE_OFN95_n429),
	.C1(n215),
	.C2(FE_OFN94_n430),
	.ZN(ALU_OPA[21]));
   OAI221_X4 U19 (.A(n417),
	.B1(FE_DBTN0_n37),
	.B2(n235),
	.C1(FE_OFN100_n391),
	.C2(n203),
	.ZN(ALU_OPB[1]));
   OAI221_X4 U20 (.A(n437),
	.B1(n66),
	.B2(n429),
	.C1(n232),
	.C2(n430),
	.ZN(ALU_OPA[4]));
   NAND3_X2 U21 (.A1(n1),
	.A2(n2),
	.A3(n3),
	.ZN(n33));
   OR3_X1 U22 (.A1(n405),
	.A2(FE_OFN23_n394),
	.A3(FE_OFN20_n393),
	.ZN(n1));
   NAND2_X1 U23 (.A1(MEM_DATA[2]),
	.A2(FE_OFN23_n394),
	.ZN(n2));
   NAND2_X1 U24 (.A1(currIMM[2]),
	.A2(FE_OFN19_n393),
	.ZN(n3));
   OAI221_X4 U28 (.A(n400),
	.B1(FE_DBTN0_n37),
	.B2(n233),
	.C1(FE_OFN100_n391),
	.C2(n202),
	.ZN(ALU_OPB[3]));
   OAI221_X2 U29 (.A(n441),
	.B1(n70),
	.B2(n429),
	.C1(n234),
	.C2(n430),
	.ZN(ALU_OPA[2]));
   OAI221_X1 U31 (.A(n402),
	.B1(FE_DBTN0_n37),
	.B2(n206),
	.C1(FE_OFN104_n391),
	.C2(n175),
	.ZN(ALU_OPB[30]));
   OAI221_X1 U32 (.A(n438),
	.B1(n68),
	.B2(n429),
	.C1(n233),
	.C2(n430),
	.ZN(ALU_OPA[3]));
   OAI221_X1 U33 (.A(n436),
	.B1(n64),
	.B2(n429),
	.C1(n231),
	.C2(n430),
	.ZN(ALU_OPA[5]));
   OAI221_X1 U34 (.A(n462),
	.B1(n54),
	.B2(n429),
	.C1(n226),
	.C2(n430),
	.ZN(ALU_OPA[10]));
   OAI221_X1 U35 (.A(n458),
	.B1(n46),
	.B2(n429),
	.C1(n222),
	.C2(n430),
	.ZN(ALU_OPA[14]));
   OAI221_X1 U36 (.A(n407),
	.B1(FE_DBTN0_n37),
	.B2(n207),
	.C1(FE_OFN104_n391),
	.C2(n176),
	.ZN(ALU_OPB[29]));
   OAI221_X1 U37 (.A(n399),
	.B1(FE_DBTN0_n37),
	.B2(n232),
	.C1(n391),
	.C2(n201),
	.ZN(ALU_OPB[4]));
   OAI221_X1 U38 (.A(n398),
	.B1(FE_DBTN0_n37),
	.B2(n231),
	.C1(n391),
	.C2(n200),
	.ZN(ALU_OPB[5]));
   OAI221_X1 U39 (.A(n397),
	.B1(FE_DBTN0_n37),
	.B2(n230),
	.C1(FE_OFN104_n391),
	.C2(n199),
	.ZN(ALU_OPB[6]));
   OAI221_X1 U40 (.A(n396),
	.B1(FE_DBTN0_n37),
	.B2(n229),
	.C1(n391),
	.C2(n198),
	.ZN(ALU_OPB[7]));
   OAI221_X1 U41 (.A(n395),
	.B1(FE_DBTN0_n37),
	.B2(n228),
	.C1(n391),
	.C2(n197),
	.ZN(ALU_OPB[8]));
   OAI221_X1 U42 (.A(n392),
	.B1(FE_DBTN0_n37),
	.B2(n227),
	.C1(n391),
	.C2(n196),
	.ZN(ALU_OPB[9]));
   OAI221_X1 U43 (.A(n427),
	.B1(FE_DBTN0_n37),
	.B2(n226),
	.C1(n391),
	.C2(n195),
	.ZN(ALU_OPB[10]));
   OAI221_X1 U44 (.A(n426),
	.B1(FE_DBTN0_n37),
	.B2(n225),
	.C1(n391),
	.C2(n194),
	.ZN(ALU_OPB[11]));
   OAI221_X1 U45 (.A(n425),
	.B1(FE_DBTN0_n37),
	.B2(n224),
	.C1(n391),
	.C2(n193),
	.ZN(ALU_OPB[12]));
   OAI221_X1 U46 (.A(n424),
	.B1(FE_DBTN0_n37),
	.B2(n223),
	.C1(FE_OFN104_n391),
	.C2(n192),
	.ZN(ALU_OPB[13]));
   OAI221_X1 U47 (.A(n423),
	.B1(FE_DBTN0_n37),
	.B2(n222),
	.C1(n391),
	.C2(n191),
	.ZN(ALU_OPB[14]));
   OAI221_X1 U48 (.A(n422),
	.B1(FE_DBTN0_n37),
	.B2(n221),
	.C1(n391),
	.C2(n190),
	.ZN(ALU_OPB[15]));
   OAI221_X1 U49 (.A(n421),
	.B1(FE_DBTN0_n37),
	.B2(n220),
	.C1(n391),
	.C2(n189),
	.ZN(ALU_OPB[16]));
   OAI221_X1 U50 (.A(n418),
	.B1(FE_DBTN0_n37),
	.B2(n217),
	.C1(FE_OFN104_n391),
	.C2(n186),
	.ZN(ALU_OPB[19]));
   OAI221_X1 U51 (.A(n416),
	.B1(FE_DBTN0_n37),
	.B2(n216),
	.C1(FE_OFN104_n391),
	.C2(n185),
	.ZN(ALU_OPB[20]));
   OAI221_X1 U52 (.A(n415),
	.B1(FE_DBTN0_n37),
	.B2(n215),
	.C1(FE_OFN104_n391),
	.C2(n184),
	.ZN(ALU_OPB[21]));
   OAI221_X1 U53 (.A(n414),
	.B1(FE_DBTN0_n37),
	.B2(n214),
	.C1(FE_OFN104_n391),
	.C2(n183),
	.ZN(ALU_OPB[22]));
   OAI221_X1 U54 (.A(n411),
	.B1(FE_DBTN0_n37),
	.B2(n211),
	.C1(FE_OFN104_n391),
	.C2(n180),
	.ZN(ALU_OPB[25]));
   OAI221_X1 U55 (.A(n410),
	.B1(FE_DBTN0_n37),
	.B2(n210),
	.C1(FE_OFN104_n391),
	.C2(n179),
	.ZN(ALU_OPB[26]));
   OAI221_X1 U56 (.A(n409),
	.B1(FE_DBTN0_n37),
	.B2(n209),
	.C1(FE_OFN104_n391),
	.C2(n178),
	.ZN(ALU_OPB[27]));
   OAI221_X1 U57 (.A(n408),
	.B1(FE_DBTN0_n37),
	.B2(n208),
	.C1(FE_OFN104_n391),
	.C2(n177),
	.ZN(ALU_OPB[28]));
   OR2_X1 U59 (.A1(n72),
	.A2(n429),
	.ZN(n5));
   OR2_X1 U60 (.A1(n235),
	.A2(n430),
	.ZN(n6));
   NAND3_X1 U61 (.A1(n5),
	.A2(n6),
	.A3(n452),
	.ZN(ALU_OPA[1]));
   AND2_X1 U62 (.A1(n172),
	.A2(n173),
	.ZN(n406));
   OR3_X1 U63 (.A1(FE_OFN19_n393),
	.A2(n8),
	.A3(n406),
	.ZN(n391));
   AND3_X1 U65 (.A1(n173),
	.A2(ALU_OPB_SEL[0]),
	.A3(ALU_OPB_SEL[1]),
	.ZN(n8));
   INV_X1 U70 (.A(n9),
	.ZN(RS2_OUT[2]));
   OAI221_X4 U86 (.A(n431),
	.B1(n56),
	.B2(n429),
	.C1(n227),
	.C2(n430),
	.ZN(ALU_OPA[9]));
   OAI221_X1 U89 (.A(n440),
	.B1(n14),
	.B2(FE_OFN95_n429),
	.C1(n206),
	.C2(FE_OFN94_n430),
	.ZN(ALU_OPA[30]));
   OAI221_X1 U90 (.A(n454),
	.B1(n38),
	.B2(FE_OFN95_n429),
	.C1(n218),
	.C2(FE_OFN94_n430),
	.ZN(ALU_OPA[18]));
   OAI221_X1 U91 (.A(n448),
	.B1(n28),
	.B2(FE_OFN95_n429),
	.C1(n213),
	.C2(FE_OFN94_n430),
	.ZN(ALU_OPA[23]));
   OAI221_X1 U92 (.A(n447),
	.B1(n26),
	.B2(FE_OFN95_n429),
	.C1(n212),
	.C2(FE_OFN94_n430),
	.ZN(ALU_OPA[24]));
   INV_X1 U118 (.A(ALU_OPA_SEL[1]),
	.ZN(n171));
   INV_X1 U123 (.A(MEM_WB_IN[4]),
	.ZN(n201));
   AOI22_X1 U124 (.A1(FE_OFN39_ALU_OPA_SEL_c_2),
	.A2(MEM_WB_IN[21]),
	.B1(FE_OFN91_n432),
	.B2(currPC[21]),
	.ZN(n450));
   AOI22_X1 U125 (.A1(FE_OFN40_ALU_OPA_SEL_c_2),
	.A2(MEM_WB_IN[20]),
	.B1(FE_OFN91_n432),
	.B2(currPC[20]),
	.ZN(n451));
   INV_X1 U126 (.A(MEM_WB_IN[18]),
	.ZN(n187));
   INV_X1 U127 (.A(MEM_WB_IN[20]),
	.ZN(n185));
   INV_X1 U128 (.A(MEM_WB_IN[16]),
	.ZN(n189));
   INV_X1 U129 (.A(MEM_WB_IN[9]),
	.ZN(n196));
   INV_X1 U130 (.A(MEM_WB_IN[19]),
	.ZN(n186));
   INV_X1 U131 (.A(EXE_MEM_IN[2]),
	.ZN(n234));
   AOI22_X1 U132 (.A1(ALU_OPA_SEL[2]),
	.A2(MEM_WB_IN[2]),
	.B1(FE_OFN90_n432),
	.B2(currPC[2]),
	.ZN(n441));
   OAI221_X1 U133 (.A(n434),
	.B1(n60),
	.B2(n429),
	.C1(n229),
	.C2(n430),
	.ZN(ALU_OPA[7]));
   OAI221_X1 U134 (.A(n433),
	.B1(n58),
	.B2(n429),
	.C1(n228),
	.C2(n430),
	.ZN(ALU_OPA[8]));
   OAI221_X1 U135 (.A(n435),
	.B1(n62),
	.B2(n429),
	.C1(n230),
	.C2(n430),
	.ZN(ALU_OPA[6]));
   INV_X1 U136 (.A(MEM_WB_IN[8]),
	.ZN(n197));
   INV_X1 U137 (.A(MEM_WB_IN[6]),
	.ZN(n199));
   INV_X1 U138 (.A(MEM_WB_IN[7]),
	.ZN(n198));
   INV_X1 U139 (.A(MEM_WB_IN[5]),
	.ZN(n200));
   OAI221_X1 U140 (.A(n420),
	.B1(FE_DBTN0_n37),
	.B2(n219),
	.C1(FE_OFN104_n391),
	.C2(n188),
	.ZN(ALU_OPB[17]));
   INV_X1 U141 (.A(MEM_WB_IN[17]),
	.ZN(n188));
   AOI221_X1 U142 (.A(n406),
	.B1(n8),
	.B2(EXE_MEM_IN[2]),
	.C1(FE_DBTN0_n37),
	.C2(MEM_WB_IN[2]),
	.ZN(n405));
   INV_X1 U143 (.A(MEM_WB_IN[3]),
	.ZN(n202));
   INV_X1 U144 (.A(MEM_WB_IN[13]),
	.ZN(n192));
   INV_X1 U145 (.A(MEM_WB_IN[14]),
	.ZN(n191));
   INV_X1 U146 (.A(MEM_WB_IN[15]),
	.ZN(n190));
   INV_X1 U147 (.A(MEM_WB_IN[0]),
	.ZN(n204));
   INV_X1 U148 (.A(MEM_WB_IN[1]),
	.ZN(n203));
   INV_X1 U149 (.A(EXE_MEM_IN[5]),
	.ZN(n231));
   INV_X1 U150 (.A(EXE_MEM_IN[3]),
	.ZN(n233));
   INV_X1 U151 (.A(EXE_MEM_IN[4]),
	.ZN(n232));
   INV_X1 U152 (.A(EXE_MEM_IN[6]),
	.ZN(n230));
   INV_X1 U153 (.A(EXE_MEM_IN[8]),
	.ZN(n228));
   INV_X1 U154 (.A(EXE_MEM_IN[7]),
	.ZN(n229));
   INV_X1 U155 (.A(EXE_MEM_IN[9]),
	.ZN(n227));
   INV_X1 U156 (.A(EXE_MEM_IN[10]),
	.ZN(n226));
   INV_X1 U157 (.A(EXE_MEM_IN[12]),
	.ZN(n224));
   INV_X1 U158 (.A(EXE_MEM_IN[14]),
	.ZN(n222));
   INV_X1 U159 (.A(EXE_MEM_IN[11]),
	.ZN(n225));
   INV_X1 U160 (.A(EXE_MEM_IN[13]),
	.ZN(n223));
   INV_X1 U161 (.A(EXE_MEM_IN[1]),
	.ZN(n235));
   INV_X1 U162 (.A(EXE_MEM_IN[0]),
	.ZN(n236));
   INV_X1 U163 (.A(MEM_WB_IN[10]),
	.ZN(n195));
   INV_X1 U164 (.A(MEM_WB_IN[12]),
	.ZN(n193));
   INV_X1 U165 (.A(MEM_WB_IN[11]),
	.ZN(n194));
   AOI22_X1 U166 (.A1(FE_OFN40_ALU_OPA_SEL_c_2),
	.A2(MEM_WB_IN[28]),
	.B1(FE_OFN91_n432),
	.B2(currPC[28]),
	.ZN(n443));
   AOI22_X1 U167 (.A1(FE_OFN39_ALU_OPA_SEL_c_2),
	.A2(MEM_WB_IN[29]),
	.B1(FE_OFN91_n432),
	.B2(currPC[29]),
	.ZN(n442));
   AOI22_X1 U168 (.A1(FE_OFN39_ALU_OPA_SEL_c_2),
	.A2(MEM_WB_IN[25]),
	.B1(FE_OFN91_n432),
	.B2(currPC[25]),
	.ZN(n446));
   AOI22_X1 U169 (.A1(FE_OFN39_ALU_OPA_SEL_c_2),
	.A2(MEM_WB_IN[27]),
	.B1(FE_OFN91_n432),
	.B2(currPC[27]),
	.ZN(n444));
   AOI22_X1 U170 (.A1(FE_OFN40_ALU_OPA_SEL_c_2),
	.A2(MEM_WB_IN[22]),
	.B1(FE_OFN91_n432),
	.B2(currPC[22]),
	.ZN(n449));
   AOI22_X1 U171 (.A1(FE_OFN39_ALU_OPA_SEL_c_2),
	.A2(MEM_WB_IN[30]),
	.B1(FE_OFN91_n432),
	.B2(currPC[30]),
	.ZN(n440));
   AOI22_X1 U172 (.A1(FE_OFN40_ALU_OPA_SEL_c_2),
	.A2(MEM_WB_IN[24]),
	.B1(FE_OFN91_n432),
	.B2(currPC[24]),
	.ZN(n447));
   AOI22_X1 U173 (.A1(FE_OFN40_ALU_OPA_SEL_c_2),
	.A2(MEM_WB_IN[26]),
	.B1(FE_OFN91_n432),
	.B2(currPC[26]),
	.ZN(n445));
   AOI22_X1 U174 (.A1(FE_OFN39_ALU_OPA_SEL_c_2),
	.A2(MEM_WB_IN[23]),
	.B1(FE_OFN91_n432),
	.B2(currPC[23]),
	.ZN(n448));
   AOI22_X1 U175 (.A1(FE_OFN39_ALU_OPA_SEL_c_2),
	.A2(MEM_WB_IN[31]),
	.B1(FE_OFN91_n432),
	.B2(currPC[31]),
	.ZN(n439));
   INV_X1 U176 (.A(MEM_WB_IN[22]),
	.ZN(n183));
   INV_X1 U177 (.A(MEM_WB_IN[26]),
	.ZN(n179));
   INV_X1 U178 (.A(MEM_WB_IN[24]),
	.ZN(n181));
   INV_X1 U179 (.A(MEM_WB_IN[21]),
	.ZN(n184));
   INV_X1 U180 (.A(MEM_WB_IN[23]),
	.ZN(n182));
   INV_X1 U181 (.A(MEM_WB_IN[25]),
	.ZN(n180));
   INV_X1 U182 (.A(MEM_WB_IN[30]),
	.ZN(n175));
   OAI221_X1 U183 (.A(n401),
	.B1(FE_DBTN0_n37),
	.B2(n205),
	.C1(FE_OFN104_n391),
	.C2(n174),
	.ZN(ALU_OPB[31]));
   INV_X1 U184 (.A(MEM_WB_IN[31]),
	.ZN(n174));
   INV_X1 U185 (.A(MEM_WB_IN[28]),
	.ZN(n177));
   INV_X1 U186 (.A(MEM_WB_IN[29]),
	.ZN(n176));
   INV_X1 U187 (.A(MEM_WB_IN[27]),
	.ZN(n178));
   INV_X1 U188 (.A(n249),
	.ZN(n529));
   AOI22_X1 U189 (.A1(RS1_IN[2]),
	.A2(FE_OFN43_n246),
	.B1(RS1_OUT[2]),
	.B2(FE_OFN0_n247),
	.ZN(n249));
   INV_X1 U190 (.A(n387),
	.ZN(n239));
   AOI22_X1 U191 (.A1(RS2_IN[2]),
	.A2(FE_OFN43_n246),
	.B1(n532),
	.B2(FE_OFN0_n247),
	.ZN(n387));
   INV_X1 U192 (.A(n245),
	.ZN(n531));
   AOI22_X1 U193 (.A1(RS1_IN[0]),
	.A2(FE_OFN43_n246),
	.B1(RS1_OUT[0]),
	.B2(FE_OFN0_n247),
	.ZN(n245));
   INV_X1 U194 (.A(n385),
	.ZN(n241));
   AOI22_X1 U195 (.A1(RS2_IN[0]),
	.A2(FE_OFN43_n246),
	.B1(RS2_OUT[0]),
	.B2(FE_OFN0_n247),
	.ZN(n385));
   INV_X1 U196 (.A(n250),
	.ZN(n528));
   AOI22_X1 U197 (.A1(RS1_IN[3]),
	.A2(FE_OFN43_n246),
	.B1(RS1_OUT[3]),
	.B2(FE_OFN0_n247),
	.ZN(n250));
   INV_X1 U198 (.A(n251),
	.ZN(n527));
   AOI22_X1 U199 (.A1(RS1_IN[4]),
	.A2(FE_OFN43_n246),
	.B1(RS1_OUT[4]),
	.B2(FE_OFN0_n247),
	.ZN(n251));
   INV_X1 U200 (.A(n304),
	.ZN(n474));
   AOI22_X1 U201 (.A1(FE_OFN2_n247),
	.A2(currPC[20]),
	.B1(FE_OFN45_n246),
	.B2(PC[20]),
	.ZN(n304));
   INV_X1 U202 (.A(n305),
	.ZN(n473));
   AOI22_X1 U203 (.A1(FE_OFN2_n247),
	.A2(currPC[21]),
	.B1(FE_OFN45_n246),
	.B2(PC[21]),
	.ZN(n305));
   INV_X1 U204 (.A(n306),
	.ZN(n472));
   AOI22_X1 U205 (.A1(FE_OFN2_n247),
	.A2(currPC[22]),
	.B1(FE_OFN45_n246),
	.B2(PC[22]),
	.ZN(n306));
   INV_X1 U206 (.A(n307),
	.ZN(n471));
   AOI22_X1 U207 (.A1(FE_OFN2_n247),
	.A2(currPC[23]),
	.B1(FE_OFN45_n246),
	.B2(PC[23]),
	.ZN(n307));
   INV_X1 U208 (.A(n308),
	.ZN(n470));
   AOI22_X1 U209 (.A1(FE_OFN2_n247),
	.A2(currPC[24]),
	.B1(FE_OFN45_n246),
	.B2(PC[24]),
	.ZN(n308));
   INV_X1 U210 (.A(n309),
	.ZN(n469));
   AOI22_X1 U211 (.A1(FE_OFN2_n247),
	.A2(currPC[25]),
	.B1(FE_OFN45_n246),
	.B2(PC[25]),
	.ZN(n309));
   INV_X1 U212 (.A(n310),
	.ZN(n468));
   AOI22_X1 U213 (.A1(FE_OFN2_n247),
	.A2(currPC[26]),
	.B1(FE_OFN45_n246),
	.B2(PC[26]),
	.ZN(n310));
   INV_X1 U214 (.A(n311),
	.ZN(n467));
   AOI22_X1 U215 (.A1(FE_OFN2_n247),
	.A2(currPC[27]),
	.B1(FE_OFN45_n246),
	.B2(PC[27]),
	.ZN(n311));
   INV_X1 U216 (.A(n312),
	.ZN(n466));
   AOI22_X1 U217 (.A1(FE_OFN2_n247),
	.A2(currPC[28]),
	.B1(FE_OFN45_n246),
	.B2(PC[28]),
	.ZN(n312));
   INV_X1 U218 (.A(n313),
	.ZN(n465));
   AOI22_X1 U219 (.A1(FE_OFN2_n247),
	.A2(currPC[29]),
	.B1(FE_OFN45_n246),
	.B2(PC[29]),
	.ZN(n313));
   INV_X1 U220 (.A(n314),
	.ZN(n464));
   AOI22_X1 U221 (.A1(FE_OFN2_n247),
	.A2(currPC[30]),
	.B1(FE_OFN45_n246),
	.B2(PC[30]),
	.ZN(n314));
   INV_X1 U222 (.A(n315),
	.ZN(n404));
   AOI22_X1 U223 (.A1(FE_OFN2_n247),
	.A2(currPC[31]),
	.B1(FE_OFN45_n246),
	.B2(PC[31]),
	.ZN(n315));
   INV_X1 U224 (.A(n388),
	.ZN(n238));
   AOI22_X1 U225 (.A1(RS2_IN[3]),
	.A2(FE_OFN43_n246),
	.B1(RS2_OUT[3]),
	.B2(FE_OFN0_n247),
	.ZN(n388));
   INV_X1 U226 (.A(n389),
	.ZN(n237));
   AOI22_X1 U227 (.A1(RS2_IN[4]),
	.A2(FE_OFN43_n246),
	.B1(RS2_OUT[4]),
	.B2(FE_OFN0_n247),
	.ZN(n389));
   NOR2_X1 U228 (.A1(en),
	.A2(rst),
	.ZN(n247));
   NOR2_X1 U229 (.A1(n247),
	.A2(rst),
	.ZN(n246));
   INV_X1 U230 (.A(EXE_MEM_IN[17]),
	.ZN(n219));
   INV_X1 U231 (.A(EXE_MEM_IN[23]),
	.ZN(n213));
   INV_X1 U232 (.A(EXE_MEM_IN[20]),
	.ZN(n216));
   INV_X1 U233 (.A(EXE_MEM_IN[21]),
	.ZN(n215));
   INV_X1 U234 (.A(EXE_MEM_IN[22]),
	.ZN(n214));
   INV_X1 U235 (.A(EXE_MEM_IN[24]),
	.ZN(n212));
   INV_X1 U236 (.A(EXE_MEM_IN[25]),
	.ZN(n211));
   INV_X1 U237 (.A(EXE_MEM_IN[15]),
	.ZN(n221));
   INV_X1 U238 (.A(EXE_MEM_IN[18]),
	.ZN(n218));
   INV_X1 U239 (.A(EXE_MEM_IN[16]),
	.ZN(n220));
   INV_X1 U240 (.A(EXE_MEM_IN[19]),
	.ZN(n217));
   INV_X1 U241 (.A(n248),
	.ZN(n530));
   AOI22_X1 U242 (.A1(RS1_IN[1]),
	.A2(FE_OFN43_n246),
	.B1(RS1_OUT[1]),
	.B2(FE_OFN0_n247),
	.ZN(n248));
   INV_X1 U243 (.A(n386),
	.ZN(n240));
   AOI22_X1 U244 (.A1(RS2_IN[1]),
	.A2(FE_OFN43_n246),
	.B1(RS2_OUT[1]),
	.B2(FE_OFN0_n247),
	.ZN(n386));
   INV_X1 U245 (.A(n373),
	.ZN(n119));
   AOI22_X1 U246 (.A1(FE_OFN2_n247),
	.A2(currRF1[25]),
	.B1(FE_OFN45_n246),
	.B2(RF_OUT1[25]),
	.ZN(n373));
   INV_X1 U247 (.A(n374),
	.ZN(n117));
   AOI22_X1 U248 (.A1(FE_OFN2_n247),
	.A2(currRF1[26]),
	.B1(FE_OFN45_n246),
	.B2(RF_OUT1[26]),
	.ZN(n374));
   INV_X1 U249 (.A(n375),
	.ZN(n115));
   AOI22_X1 U250 (.A1(FE_OFN2_n247),
	.A2(currRF1[27]),
	.B1(FE_OFN45_n246),
	.B2(RF_OUT1[27]),
	.ZN(n375));
   INV_X1 U251 (.A(n376),
	.ZN(n113));
   AOI22_X1 U252 (.A1(FE_OFN2_n247),
	.A2(currRF1[28]),
	.B1(FE_OFN45_n246),
	.B2(RF_OUT1[28]),
	.ZN(n376));
   INV_X1 U253 (.A(n377),
	.ZN(n111));
   AOI22_X1 U254 (.A1(FE_OFN2_n247),
	.A2(currRF1[29]),
	.B1(FE_OFN45_n246),
	.B2(RF_OUT1[29]),
	.ZN(n377));
   INV_X1 U255 (.A(n378),
	.ZN(n109));
   AOI22_X1 U256 (.A1(FE_OFN2_n247),
	.A2(currRF1[30]),
	.B1(FE_OFN45_n246),
	.B2(RF_OUT1[30]),
	.ZN(n378));
   INV_X1 U257 (.A(n380),
	.ZN(n403));
   AOI22_X1 U258 (.A1(RD_IN[0]),
	.A2(FE_OFN43_n246),
	.B1(RD_OUT[0]),
	.B2(n247),
	.ZN(n380));
   INV_X1 U259 (.A(n381),
	.ZN(n390));
   AOI22_X1 U260 (.A1(RD_IN[1]),
	.A2(FE_OFN43_n246),
	.B1(RD_OUT[1]),
	.B2(FE_OFN0_n247),
	.ZN(n381));
   INV_X1 U261 (.A(n382),
	.ZN(n244));
   AOI22_X1 U262 (.A1(RD_IN[2]),
	.A2(FE_OFN43_n246),
	.B1(RD_OUT[2]),
	.B2(n247),
	.ZN(n382));
   INV_X1 U263 (.A(n283),
	.ZN(n495));
   AOI22_X1 U264 (.A1(FE_OFN2_n247),
	.A2(currIMM[31]),
	.B1(FE_OFN45_n246),
	.B2(IMM[31]),
	.ZN(n283));
   INV_X1 U265 (.A(n252),
	.ZN(n526));
   AOI22_X1 U266 (.A1(FE_OFN0_n247),
	.A2(currIMM[0]),
	.B1(FE_OFN43_n246),
	.B2(IMM[0]),
	.ZN(n252));
   INV_X1 U267 (.A(n383),
	.ZN(n243));
   AOI22_X1 U268 (.A1(RD_IN[3]),
	.A2(FE_OFN43_n246),
	.B1(RD_OUT[3]),
	.B2(FE_OFN0_n247),
	.ZN(n383));
   INV_X1 U269 (.A(n384),
	.ZN(n242));
   AOI22_X1 U270 (.A1(RD_IN[4]),
	.A2(FE_OFN43_n246),
	.B1(RD_OUT[4]),
	.B2(n247),
	.ZN(n384));
   INV_X1 U271 (.A(n281),
	.ZN(n497));
   AOI22_X1 U272 (.A1(FE_OFN2_n247),
	.A2(currIMM[29]),
	.B1(FE_OFN45_n246),
	.B2(IMM[29]),
	.ZN(n281));
   INV_X1 U273 (.A(n316),
	.ZN(n170));
   AOI22_X1 U274 (.A1(FE_OFN1_n247),
	.A2(MEM_DATA[0]),
	.B1(FE_OFN44_n246),
	.B2(RF_OUT2[0]),
	.ZN(n316));
   INV_X1 U275 (.A(n317),
	.ZN(n168));
   AOI22_X1 U276 (.A1(FE_OFN2_n247),
	.A2(MEM_DATA[1]),
	.B1(FE_OFN45_n246),
	.B2(RF_OUT2[1]),
	.ZN(n317));
   INV_X1 U277 (.A(n318),
	.ZN(n166));
   AOI22_X1 U278 (.A1(FE_OFN2_n247),
	.A2(MEM_DATA[2]),
	.B1(FE_OFN45_n246),
	.B2(RF_OUT2[2]),
	.ZN(n318));
   INV_X1 U279 (.A(n319),
	.ZN(n164));
   AOI22_X1 U280 (.A1(FE_OFN1_n247),
	.A2(MEM_DATA[3]),
	.B1(FE_OFN44_n246),
	.B2(RF_OUT2[3]),
	.ZN(n319));
   INV_X1 U281 (.A(n320),
	.ZN(n162));
   AOI22_X1 U282 (.A1(FE_OFN0_n247),
	.A2(MEM_DATA[4]),
	.B1(FE_OFN43_n246),
	.B2(RF_OUT2[4]),
	.ZN(n320));
   INV_X1 U283 (.A(n321),
	.ZN(n160));
   AOI22_X1 U284 (.A1(FE_OFN1_n247),
	.A2(MEM_DATA[5]),
	.B1(FE_OFN44_n246),
	.B2(RF_OUT2[5]),
	.ZN(n321));
   INV_X1 U285 (.A(n322),
	.ZN(n158));
   AOI22_X1 U286 (.A1(FE_OFN1_n247),
	.A2(MEM_DATA[6]),
	.B1(FE_OFN44_n246),
	.B2(RF_OUT2[6]),
	.ZN(n322));
   INV_X1 U287 (.A(n323),
	.ZN(n156));
   AOI22_X1 U288 (.A1(FE_OFN1_n247),
	.A2(MEM_DATA[7]),
	.B1(FE_OFN44_n246),
	.B2(RF_OUT2[7]),
	.ZN(n323));
   INV_X1 U289 (.A(n324),
	.ZN(n154));
   AOI22_X1 U290 (.A1(FE_OFN1_n247),
	.A2(MEM_DATA[8]),
	.B1(FE_OFN44_n246),
	.B2(RF_OUT2[8]),
	.ZN(n324));
   INV_X1 U291 (.A(n325),
	.ZN(n152));
   AOI22_X1 U292 (.A1(FE_OFN1_n247),
	.A2(MEM_DATA[9]),
	.B1(FE_OFN44_n246),
	.B2(RF_OUT2[9]),
	.ZN(n325));
   INV_X1 U293 (.A(n326),
	.ZN(n150));
   AOI22_X1 U294 (.A1(FE_OFN1_n247),
	.A2(MEM_DATA[10]),
	.B1(FE_OFN44_n246),
	.B2(RF_OUT2[10]),
	.ZN(n326));
   INV_X1 U295 (.A(n327),
	.ZN(n148));
   AOI22_X1 U296 (.A1(FE_OFN0_n247),
	.A2(MEM_DATA[11]),
	.B1(FE_OFN43_n246),
	.B2(RF_OUT2[11]),
	.ZN(n327));
   INV_X1 U297 (.A(n328),
	.ZN(n146));
   AOI22_X1 U298 (.A1(FE_OFN1_n247),
	.A2(MEM_DATA[12]),
	.B1(FE_OFN44_n246),
	.B2(RF_OUT2[12]),
	.ZN(n328));
   INV_X1 U299 (.A(n329),
	.ZN(n144));
   AOI22_X1 U300 (.A1(FE_OFN1_n247),
	.A2(MEM_DATA[13]),
	.B1(FE_OFN44_n246),
	.B2(RF_OUT2[13]),
	.ZN(n329));
   INV_X1 U301 (.A(n330),
	.ZN(n142));
   AOI22_X1 U302 (.A1(FE_OFN0_n247),
	.A2(MEM_DATA[14]),
	.B1(FE_OFN43_n246),
	.B2(RF_OUT2[14]),
	.ZN(n330));
   INV_X1 U303 (.A(n331),
	.ZN(n140));
   AOI22_X1 U304 (.A1(FE_OFN0_n247),
	.A2(MEM_DATA[15]),
	.B1(FE_OFN43_n246),
	.B2(RF_OUT2[15]),
	.ZN(n331));
   INV_X1 U305 (.A(n332),
	.ZN(n138));
   AOI22_X1 U306 (.A1(FE_OFN1_n247),
	.A2(MEM_DATA[16]),
	.B1(FE_OFN44_n246),
	.B2(RF_OUT2[16]),
	.ZN(n332));
   INV_X1 U307 (.A(n333),
	.ZN(n136));
   AOI22_X1 U308 (.A1(FE_OFN2_n247),
	.A2(MEM_DATA[17]),
	.B1(FE_OFN45_n246),
	.B2(RF_OUT2[17]),
	.ZN(n333));
   INV_X1 U309 (.A(n334),
	.ZN(n134));
   AOI22_X1 U310 (.A1(FE_OFN2_n247),
	.A2(MEM_DATA[18]),
	.B1(FE_OFN45_n246),
	.B2(RF_OUT2[18]),
	.ZN(n334));
   INV_X1 U311 (.A(n335),
	.ZN(n132));
   AOI22_X1 U312 (.A1(FE_OFN2_n247),
	.A2(MEM_DATA[19]),
	.B1(FE_OFN45_n246),
	.B2(RF_OUT2[19]),
	.ZN(n335));
   INV_X1 U313 (.A(n336),
	.ZN(n130));
   AOI22_X1 U314 (.A1(FE_OFN2_n247),
	.A2(MEM_DATA[20]),
	.B1(FE_OFN45_n246),
	.B2(RF_OUT2[20]),
	.ZN(n336));
   INV_X1 U315 (.A(n337),
	.ZN(n128));
   AOI22_X1 U316 (.A1(FE_OFN2_n247),
	.A2(MEM_DATA[21]),
	.B1(FE_OFN45_n246),
	.B2(RF_OUT2[21]),
	.ZN(n337));
   INV_X1 U317 (.A(n338),
	.ZN(n126));
   AOI22_X1 U318 (.A1(FE_OFN2_n247),
	.A2(MEM_DATA[22]),
	.B1(FE_OFN45_n246),
	.B2(RF_OUT2[22]),
	.ZN(n338));
   INV_X1 U319 (.A(n339),
	.ZN(n124));
   AOI22_X1 U320 (.A1(FE_OFN2_n247),
	.A2(MEM_DATA[23]),
	.B1(FE_OFN45_n246),
	.B2(RF_OUT2[23]),
	.ZN(n339));
   INV_X1 U321 (.A(n340),
	.ZN(n122));
   AOI22_X1 U322 (.A1(FE_OFN2_n247),
	.A2(MEM_DATA[24]),
	.B1(FE_OFN45_n246),
	.B2(RF_OUT2[24]),
	.ZN(n340));
   INV_X1 U323 (.A(n341),
	.ZN(n120));
   AOI22_X1 U324 (.A1(FE_OFN2_n247),
	.A2(MEM_DATA[25]),
	.B1(FE_OFN45_n246),
	.B2(RF_OUT2[25]),
	.ZN(n341));
   INV_X1 U325 (.A(n342),
	.ZN(n118));
   AOI22_X1 U326 (.A1(FE_OFN2_n247),
	.A2(MEM_DATA[26]),
	.B1(FE_OFN45_n246),
	.B2(RF_OUT2[26]),
	.ZN(n342));
   INV_X1 U327 (.A(n343),
	.ZN(n116));
   AOI22_X1 U328 (.A1(FE_OFN2_n247),
	.A2(MEM_DATA[27]),
	.B1(FE_OFN45_n246),
	.B2(RF_OUT2[27]),
	.ZN(n343));
   INV_X1 U329 (.A(n344),
	.ZN(n114));
   AOI22_X1 U330 (.A1(FE_OFN2_n247),
	.A2(MEM_DATA[28]),
	.B1(FE_OFN45_n246),
	.B2(RF_OUT2[28]),
	.ZN(n344));
   INV_X1 U331 (.A(n345),
	.ZN(n112));
   AOI22_X1 U332 (.A1(FE_OFN2_n247),
	.A2(MEM_DATA[29]),
	.B1(FE_OFN45_n246),
	.B2(RF_OUT2[29]),
	.ZN(n345));
   INV_X1 U333 (.A(n346),
	.ZN(n110));
   AOI22_X1 U334 (.A1(FE_OFN2_n247),
	.A2(MEM_DATA[30]),
	.B1(FE_OFN45_n246),
	.B2(RF_OUT2[30]),
	.ZN(n346));
   INV_X1 U335 (.A(n347),
	.ZN(n108));
   AOI22_X1 U336 (.A1(FE_OFN2_n247),
	.A2(MEM_DATA[31]),
	.B1(FE_OFN45_n246),
	.B2(RF_OUT2[31]),
	.ZN(n347));
   INV_X1 U337 (.A(n348),
	.ZN(n169));
   AOI22_X1 U338 (.A1(FE_OFN1_n247),
	.A2(currRF1[0]),
	.B1(FE_OFN44_n246),
	.B2(RF_OUT1[0]),
	.ZN(n348));
   INV_X1 U339 (.A(n349),
	.ZN(n167));
   AOI22_X1 U340 (.A1(FE_OFN2_n247),
	.A2(currRF1[1]),
	.B1(FE_OFN45_n246),
	.B2(RF_OUT1[1]),
	.ZN(n349));
   INV_X1 U341 (.A(n350),
	.ZN(n165));
   AOI22_X1 U342 (.A1(FE_OFN2_n247),
	.A2(currRF1[2]),
	.B1(FE_OFN45_n246),
	.B2(RF_OUT1[2]),
	.ZN(n350));
   INV_X1 U343 (.A(n351),
	.ZN(n163));
   AOI22_X1 U344 (.A1(FE_OFN1_n247),
	.A2(currRF1[3]),
	.B1(FE_OFN44_n246),
	.B2(RF_OUT1[3]),
	.ZN(n351));
   INV_X1 U345 (.A(n352),
	.ZN(n161));
   AOI22_X1 U346 (.A1(FE_OFN0_n247),
	.A2(currRF1[4]),
	.B1(FE_OFN43_n246),
	.B2(RF_OUT1[4]),
	.ZN(n352));
   INV_X1 U347 (.A(n353),
	.ZN(n159));
   AOI22_X1 U348 (.A1(FE_OFN1_n247),
	.A2(currRF1[5]),
	.B1(FE_OFN44_n246),
	.B2(RF_OUT1[5]),
	.ZN(n353));
   INV_X1 U349 (.A(n354),
	.ZN(n157));
   AOI22_X1 U350 (.A1(FE_OFN1_n247),
	.A2(currRF1[6]),
	.B1(FE_OFN44_n246),
	.B2(RF_OUT1[6]),
	.ZN(n354));
   INV_X1 U351 (.A(n355),
	.ZN(n155));
   AOI22_X1 U352 (.A1(FE_OFN1_n247),
	.A2(currRF1[7]),
	.B1(FE_OFN44_n246),
	.B2(RF_OUT1[7]),
	.ZN(n355));
   INV_X1 U353 (.A(n356),
	.ZN(n153));
   AOI22_X1 U354 (.A1(FE_OFN1_n247),
	.A2(currRF1[8]),
	.B1(FE_OFN44_n246),
	.B2(RF_OUT1[8]),
	.ZN(n356));
   INV_X1 U355 (.A(n357),
	.ZN(n151));
   AOI22_X1 U356 (.A1(FE_OFN1_n247),
	.A2(currRF1[9]),
	.B1(FE_OFN44_n246),
	.B2(RF_OUT1[9]),
	.ZN(n357));
   INV_X1 U357 (.A(n358),
	.ZN(n149));
   AOI22_X1 U358 (.A1(FE_OFN1_n247),
	.A2(currRF1[10]),
	.B1(FE_OFN44_n246),
	.B2(RF_OUT1[10]),
	.ZN(n358));
   INV_X1 U359 (.A(n359),
	.ZN(n147));
   AOI22_X1 U360 (.A1(FE_OFN0_n247),
	.A2(currRF1[11]),
	.B1(FE_OFN44_n246),
	.B2(RF_OUT1[11]),
	.ZN(n359));
   INV_X1 U361 (.A(n360),
	.ZN(n145));
   AOI22_X1 U362 (.A1(FE_OFN1_n247),
	.A2(currRF1[12]),
	.B1(FE_OFN44_n246),
	.B2(RF_OUT1[12]),
	.ZN(n360));
   INV_X1 U363 (.A(n361),
	.ZN(n143));
   AOI22_X1 U364 (.A1(FE_OFN1_n247),
	.A2(currRF1[13]),
	.B1(FE_OFN45_n246),
	.B2(RF_OUT1[13]),
	.ZN(n361));
   INV_X1 U365 (.A(n362),
	.ZN(n141));
   AOI22_X1 U366 (.A1(FE_OFN0_n247),
	.A2(currRF1[14]),
	.B1(FE_OFN43_n246),
	.B2(RF_OUT1[14]),
	.ZN(n362));
   INV_X1 U367 (.A(n363),
	.ZN(n139));
   AOI22_X1 U368 (.A1(FE_OFN0_n247),
	.A2(currRF1[15]),
	.B1(FE_OFN44_n246),
	.B2(RF_OUT1[15]),
	.ZN(n363));
   INV_X1 U369 (.A(n364),
	.ZN(n137));
   AOI22_X1 U370 (.A1(FE_OFN1_n247),
	.A2(currRF1[16]),
	.B1(FE_OFN44_n246),
	.B2(RF_OUT1[16]),
	.ZN(n364));
   INV_X1 U371 (.A(n365),
	.ZN(n135));
   AOI22_X1 U372 (.A1(FE_OFN2_n247),
	.A2(currRF1[17]),
	.B1(FE_OFN45_n246),
	.B2(RF_OUT1[17]),
	.ZN(n365));
   INV_X1 U373 (.A(n366),
	.ZN(n133));
   AOI22_X1 U374 (.A1(FE_OFN2_n247),
	.A2(currRF1[18]),
	.B1(FE_OFN45_n246),
	.B2(RF_OUT1[18]),
	.ZN(n366));
   INV_X1 U375 (.A(n367),
	.ZN(n131));
   AOI22_X1 U376 (.A1(FE_OFN2_n247),
	.A2(currRF1[19]),
	.B1(FE_OFN45_n246),
	.B2(RF_OUT1[19]),
	.ZN(n367));
   INV_X1 U377 (.A(n368),
	.ZN(n129));
   AOI22_X1 U378 (.A1(FE_OFN2_n247),
	.A2(currRF1[20]),
	.B1(FE_OFN45_n246),
	.B2(RF_OUT1[20]),
	.ZN(n368));
   INV_X1 U379 (.A(n369),
	.ZN(n127));
   AOI22_X1 U380 (.A1(FE_OFN2_n247),
	.A2(currRF1[21]),
	.B1(FE_OFN45_n246),
	.B2(RF_OUT1[21]),
	.ZN(n369));
   INV_X1 U381 (.A(n370),
	.ZN(n125));
   AOI22_X1 U382 (.A1(FE_OFN2_n247),
	.A2(currRF1[22]),
	.B1(FE_OFN45_n246),
	.B2(RF_OUT1[22]),
	.ZN(n370));
   INV_X1 U383 (.A(n371),
	.ZN(n123));
   AOI22_X1 U384 (.A1(FE_OFN2_n247),
	.A2(currRF1[23]),
	.B1(FE_OFN45_n246),
	.B2(RF_OUT1[23]),
	.ZN(n371));
   INV_X1 U385 (.A(n372),
	.ZN(n121));
   AOI22_X1 U386 (.A1(FE_OFN2_n247),
	.A2(currRF1[24]),
	.B1(FE_OFN45_n246),
	.B2(RF_OUT1[24]),
	.ZN(n372));
   INV_X1 U387 (.A(n261),
	.ZN(n517));
   AOI22_X1 U388 (.A1(FE_OFN0_n247),
	.A2(currIMM[9]),
	.B1(FE_OFN43_n246),
	.B2(IMM[9]),
	.ZN(n261));
   INV_X1 U389 (.A(n262),
	.ZN(n516));
   AOI22_X1 U390 (.A1(FE_OFN0_n247),
	.A2(currIMM[10]),
	.B1(FE_OFN43_n246),
	.B2(IMM[10]),
	.ZN(n262));
   INV_X1 U391 (.A(n263),
	.ZN(n515));
   AOI22_X1 U392 (.A1(FE_OFN0_n247),
	.A2(currIMM[11]),
	.B1(FE_OFN43_n246),
	.B2(IMM[11]),
	.ZN(n263));
   INV_X1 U393 (.A(n264),
	.ZN(n514));
   AOI22_X1 U394 (.A1(FE_OFN0_n247),
	.A2(currIMM[12]),
	.B1(FE_OFN43_n246),
	.B2(IMM[12]),
	.ZN(n264));
   INV_X1 U395 (.A(n265),
	.ZN(n513));
   AOI22_X1 U396 (.A1(FE_OFN0_n247),
	.A2(currIMM[13]),
	.B1(FE_OFN43_n246),
	.B2(IMM[13]),
	.ZN(n265));
   INV_X1 U397 (.A(n266),
	.ZN(n512));
   AOI22_X1 U398 (.A1(FE_OFN0_n247),
	.A2(currIMM[14]),
	.B1(FE_OFN43_n246),
	.B2(IMM[14]),
	.ZN(n266));
   INV_X1 U399 (.A(n267),
	.ZN(n511));
   AOI22_X1 U400 (.A1(FE_OFN0_n247),
	.A2(currIMM[15]),
	.B1(FE_OFN43_n246),
	.B2(IMM[15]),
	.ZN(n267));
   INV_X1 U401 (.A(n268),
	.ZN(n510));
   AOI22_X1 U402 (.A1(FE_OFN0_n247),
	.A2(currIMM[16]),
	.B1(FE_OFN43_n246),
	.B2(IMM[16]),
	.ZN(n268));
   INV_X1 U403 (.A(n269),
	.ZN(n509));
   AOI22_X1 U404 (.A1(FE_OFN0_n247),
	.A2(currIMM[17]),
	.B1(FE_OFN43_n246),
	.B2(IMM[17]),
	.ZN(n269));
   INV_X1 U405 (.A(n270),
	.ZN(n508));
   AOI22_X1 U406 (.A1(FE_OFN0_n247),
	.A2(currIMM[18]),
	.B1(FE_OFN43_n246),
	.B2(IMM[18]),
	.ZN(n270));
   INV_X1 U407 (.A(n271),
	.ZN(n507));
   AOI22_X1 U408 (.A1(FE_OFN2_n247),
	.A2(currIMM[19]),
	.B1(FE_OFN45_n246),
	.B2(IMM[19]),
	.ZN(n271));
   INV_X1 U409 (.A(n272),
	.ZN(n506));
   AOI22_X1 U410 (.A1(FE_OFN2_n247),
	.A2(currIMM[20]),
	.B1(FE_OFN45_n246),
	.B2(IMM[20]),
	.ZN(n272));
   INV_X1 U411 (.A(n273),
	.ZN(n505));
   AOI22_X1 U412 (.A1(FE_OFN2_n247),
	.A2(currIMM[21]),
	.B1(FE_OFN45_n246),
	.B2(IMM[21]),
	.ZN(n273));
   INV_X1 U413 (.A(n274),
	.ZN(n504));
   AOI22_X1 U414 (.A1(FE_OFN2_n247),
	.A2(currIMM[22]),
	.B1(FE_OFN45_n246),
	.B2(IMM[22]),
	.ZN(n274));
   INV_X1 U415 (.A(n275),
	.ZN(n503));
   AOI22_X1 U416 (.A1(FE_OFN2_n247),
	.A2(currIMM[23]),
	.B1(FE_OFN45_n246),
	.B2(IMM[23]),
	.ZN(n275));
   INV_X1 U417 (.A(n276),
	.ZN(n502));
   AOI22_X1 U418 (.A1(FE_OFN2_n247),
	.A2(currIMM[24]),
	.B1(FE_OFN45_n246),
	.B2(IMM[24]),
	.ZN(n276));
   INV_X1 U419 (.A(n277),
	.ZN(n501));
   AOI22_X1 U420 (.A1(FE_OFN2_n247),
	.A2(currIMM[25]),
	.B1(FE_OFN45_n246),
	.B2(IMM[25]),
	.ZN(n277));
   INV_X1 U421 (.A(n278),
	.ZN(n500));
   AOI22_X1 U422 (.A1(FE_OFN2_n247),
	.A2(currIMM[26]),
	.B1(FE_OFN45_n246),
	.B2(IMM[26]),
	.ZN(n278));
   INV_X1 U423 (.A(n279),
	.ZN(n499));
   AOI22_X1 U424 (.A1(FE_OFN2_n247),
	.A2(currIMM[27]),
	.B1(FE_OFN45_n246),
	.B2(IMM[27]),
	.ZN(n279));
   INV_X1 U425 (.A(n280),
	.ZN(n498));
   AOI22_X1 U426 (.A1(FE_OFN2_n247),
	.A2(currIMM[28]),
	.B1(FE_OFN45_n246),
	.B2(IMM[28]),
	.ZN(n280));
   INV_X1 U427 (.A(n282),
	.ZN(n496));
   AOI22_X1 U428 (.A1(FE_OFN2_n247),
	.A2(currIMM[30]),
	.B1(FE_OFN45_n246),
	.B2(IMM[30]),
	.ZN(n282));
   INV_X1 U429 (.A(n284),
	.ZN(n494));
   AOI22_X1 U430 (.A1(FE_OFN0_n247),
	.A2(currPC[0]),
	.B1(FE_OFN43_n246),
	.B2(PC[0]),
	.ZN(n284));
   INV_X1 U431 (.A(n285),
	.ZN(n493));
   AOI22_X1 U432 (.A1(FE_OFN0_n247),
	.A2(currPC[1]),
	.B1(FE_OFN43_n246),
	.B2(PC[1]),
	.ZN(n285));
   INV_X1 U433 (.A(n286),
	.ZN(n492));
   AOI22_X1 U434 (.A1(FE_OFN0_n247),
	.A2(currPC[2]),
	.B1(FE_OFN43_n246),
	.B2(PC[2]),
	.ZN(n286));
   INV_X1 U435 (.A(n287),
	.ZN(n491));
   AOI22_X1 U436 (.A1(FE_OFN0_n247),
	.A2(currPC[3]),
	.B1(FE_OFN43_n246),
	.B2(PC[3]),
	.ZN(n287));
   INV_X1 U437 (.A(n288),
	.ZN(n490));
   AOI22_X1 U438 (.A1(FE_OFN0_n247),
	.A2(currPC[4]),
	.B1(FE_OFN43_n246),
	.B2(PC[4]),
	.ZN(n288));
   INV_X1 U439 (.A(n289),
	.ZN(n489));
   AOI22_X1 U440 (.A1(FE_OFN0_n247),
	.A2(currPC[5]),
	.B1(FE_OFN43_n246),
	.B2(PC[5]),
	.ZN(n289));
   INV_X1 U441 (.A(n290),
	.ZN(n488));
   AOI22_X1 U442 (.A1(FE_OFN0_n247),
	.A2(currPC[6]),
	.B1(FE_OFN43_n246),
	.B2(PC[6]),
	.ZN(n290));
   INV_X1 U443 (.A(n291),
	.ZN(n487));
   AOI22_X1 U444 (.A1(FE_OFN0_n247),
	.A2(currPC[7]),
	.B1(FE_OFN43_n246),
	.B2(PC[7]),
	.ZN(n291));
   INV_X1 U445 (.A(n292),
	.ZN(n486));
   AOI22_X1 U446 (.A1(FE_OFN0_n247),
	.A2(currPC[8]),
	.B1(FE_OFN43_n246),
	.B2(PC[8]),
	.ZN(n292));
   INV_X1 U447 (.A(n293),
	.ZN(n485));
   AOI22_X1 U448 (.A1(FE_OFN0_n247),
	.A2(currPC[9]),
	.B1(FE_OFN43_n246),
	.B2(PC[9]),
	.ZN(n293));
   INV_X1 U449 (.A(n294),
	.ZN(n484));
   AOI22_X1 U450 (.A1(FE_OFN0_n247),
	.A2(currPC[10]),
	.B1(FE_OFN43_n246),
	.B2(PC[10]),
	.ZN(n294));
   INV_X1 U451 (.A(n295),
	.ZN(n483));
   AOI22_X1 U452 (.A1(FE_OFN0_n247),
	.A2(currPC[11]),
	.B1(FE_OFN43_n246),
	.B2(PC[11]),
	.ZN(n295));
   INV_X1 U453 (.A(n296),
	.ZN(n482));
   AOI22_X1 U454 (.A1(FE_OFN0_n247),
	.A2(currPC[12]),
	.B1(FE_OFN43_n246),
	.B2(PC[12]),
	.ZN(n296));
   INV_X1 U455 (.A(n297),
	.ZN(n481));
   AOI22_X1 U456 (.A1(FE_OFN0_n247),
	.A2(currPC[13]),
	.B1(FE_OFN43_n246),
	.B2(PC[13]),
	.ZN(n297));
   INV_X1 U457 (.A(n298),
	.ZN(n480));
   AOI22_X1 U458 (.A1(FE_OFN0_n247),
	.A2(currPC[14]),
	.B1(FE_OFN43_n246),
	.B2(PC[14]),
	.ZN(n298));
   INV_X1 U459 (.A(n299),
	.ZN(n479));
   AOI22_X1 U460 (.A1(FE_OFN0_n247),
	.A2(currPC[15]),
	.B1(FE_OFN43_n246),
	.B2(PC[15]),
	.ZN(n299));
   INV_X1 U461 (.A(n300),
	.ZN(n478));
   AOI22_X1 U462 (.A1(FE_OFN0_n247),
	.A2(currPC[16]),
	.B1(FE_OFN43_n246),
	.B2(PC[16]),
	.ZN(n300));
   INV_X1 U463 (.A(n301),
	.ZN(n477));
   AOI22_X1 U464 (.A1(FE_OFN0_n247),
	.A2(currPC[17]),
	.B1(FE_OFN43_n246),
	.B2(PC[17]),
	.ZN(n301));
   INV_X1 U465 (.A(n302),
	.ZN(n476));
   AOI22_X1 U466 (.A1(FE_OFN2_n247),
	.A2(currPC[18]),
	.B1(FE_OFN45_n246),
	.B2(PC[18]),
	.ZN(n302));
   INV_X1 U467 (.A(n303),
	.ZN(n475));
   AOI22_X1 U468 (.A1(FE_OFN2_n247),
	.A2(currPC[19]),
	.B1(FE_OFN45_n246),
	.B2(PC[19]),
	.ZN(n303));
   INV_X1 U469 (.A(n253),
	.ZN(n525));
   AOI22_X1 U470 (.A1(FE_OFN0_n247),
	.A2(currIMM[1]),
	.B1(FE_OFN43_n246),
	.B2(IMM[1]),
	.ZN(n253));
   INV_X1 U471 (.A(n254),
	.ZN(n524));
   AOI22_X1 U472 (.A1(FE_OFN0_n247),
	.A2(currIMM[2]),
	.B1(FE_OFN43_n246),
	.B2(IMM[2]),
	.ZN(n254));
   INV_X1 U473 (.A(n255),
	.ZN(n523));
   AOI22_X1 U474 (.A1(FE_OFN0_n247),
	.A2(currIMM[3]),
	.B1(FE_OFN43_n246),
	.B2(IMM[3]),
	.ZN(n255));
   INV_X1 U475 (.A(n256),
	.ZN(n522));
   AOI22_X1 U476 (.A1(FE_OFN0_n247),
	.A2(currIMM[4]),
	.B1(FE_OFN43_n246),
	.B2(IMM[4]),
	.ZN(n256));
   INV_X1 U477 (.A(n257),
	.ZN(n521));
   AOI22_X1 U478 (.A1(FE_OFN0_n247),
	.A2(currIMM[5]),
	.B1(FE_OFN43_n246),
	.B2(IMM[5]),
	.ZN(n257));
   INV_X1 U479 (.A(n258),
	.ZN(n520));
   AOI22_X1 U480 (.A1(FE_OFN0_n247),
	.A2(currIMM[6]),
	.B1(FE_OFN43_n246),
	.B2(IMM[6]),
	.ZN(n258));
   INV_X1 U481 (.A(n259),
	.ZN(n519));
   AOI22_X1 U482 (.A1(FE_OFN0_n247),
	.A2(currIMM[7]),
	.B1(FE_OFN43_n246),
	.B2(IMM[7]),
	.ZN(n259));
   INV_X1 U483 (.A(n260),
	.ZN(n518));
   AOI22_X1 U484 (.A1(FE_OFN0_n247),
	.A2(currIMM[8]),
	.B1(FE_OFN43_n246),
	.B2(IMM[8]),
	.ZN(n260));
   INV_X1 U485 (.A(n379),
	.ZN(n107));
   AOI22_X1 U486 (.A1(FE_OFN2_n247),
	.A2(currRF1[31]),
	.B1(FE_OFN45_n246),
	.B2(RF_OUT1[31]),
	.ZN(n379));
   INV_X1 U487 (.A(EXE_MEM_IN[30]),
	.ZN(n206));
   INV_X1 U488 (.A(EXE_MEM_IN[28]),
	.ZN(n208));
   INV_X1 U489 (.A(EXE_MEM_IN[27]),
	.ZN(n209));
   INV_X1 U490 (.A(EXE_MEM_IN[29]),
	.ZN(n207));
   INV_X1 U491 (.A(EXE_MEM_IN[31]),
	.ZN(n205));
   INV_X1 U492 (.A(EXE_MEM_IN[26]),
	.ZN(n210));
   AOI22_X1 U493 (.A1(ALU_OPA_SEL[2]),
	.A2(MEM_WB_IN[9]),
	.B1(FE_OFN90_n432),
	.B2(currPC[9]),
	.ZN(n431));
   AOI22_X1 U494 (.A1(ALU_OPA_SEL[2]),
	.A2(MEM_WB_IN[8]),
	.B1(FE_OFN90_n432),
	.B2(currPC[8]),
	.ZN(n433));
   AOI22_X1 U497 (.A1(ALU_OPA_SEL[2]),
	.A2(MEM_WB_IN[7]),
	.B1(FE_OFN90_n432),
	.B2(currPC[7]),
	.ZN(n434));
   AOI22_X1 U498 (.A1(FE_OFN39_ALU_OPA_SEL_c_2),
	.A2(MEM_WB_IN[6]),
	.B1(FE_OFN90_n432),
	.B2(currPC[6]),
	.ZN(n435));
   AOI22_X1 U499 (.A1(ALU_OPA_SEL[2]),
	.A2(MEM_WB_IN[5]),
	.B1(FE_OFN90_n432),
	.B2(currPC[5]),
	.ZN(n436));
   AOI22_X1 U500 (.A1(ALU_OPA_SEL[2]),
	.A2(MEM_WB_IN[4]),
	.B1(FE_OFN90_n432),
	.B2(currPC[4]),
	.ZN(n437));
   AOI22_X1 U501 (.A1(ALU_OPA_SEL[2]),
	.A2(MEM_WB_IN[3]),
	.B1(FE_OFN90_n432),
	.B2(currPC[3]),
	.ZN(n438));
   INV_X1 U502 (.A(ALU_OPB_SEL[2]),
	.ZN(n173));
   OAI221_X1 U505 (.A(n460),
	.B1(n50),
	.B2(n429),
	.C1(n224),
	.C2(n430),
	.ZN(ALU_OPA[12]));
   OAI221_X1 U507 (.A(n412),
	.B1(FE_DBTN0_n37),
	.B2(n212),
	.C1(FE_OFN104_n391),
	.C2(n181),
	.ZN(ALU_OPB[24]));
   OAI221_X1 U508 (.A(n413),
	.B1(FE_DBTN0_n37),
	.B2(n213),
	.C1(FE_OFN104_n391),
	.C2(n182),
	.ZN(ALU_OPB[23]));
   OAI221_X1 U509 (.A(n419),
	.B1(FE_DBTN0_n37),
	.B2(n218),
	.C1(FE_OFN104_n391),
	.C2(n187),
	.ZN(ALU_OPB[18]));
   NOR3_X1 U511 (.A1(n172),
	.A2(ALU_OPB_SEL[2]),
	.A3(ALU_OPB_SEL[1]),
	.ZN(n393));
   NOR3_X1 U512 (.A1(ALU_OPA_SEL[1]),
	.A2(ALU_OPA_SEL[0]),
	.A3(ALU_OPA_SEL[2]),
	.ZN(n55));
   AOI22_X1 U514 (.A1(FE_OFN20_n393),
	.A2(currIMM[17]),
	.B1(FE_OFN28_n394),
	.B2(MEM_DATA[17]),
	.ZN(n420));
   AOI22_X1 U515 (.A1(FE_OFN20_n393),
	.A2(currIMM[13]),
	.B1(FE_OFN23_n394),
	.B2(MEM_DATA[13]),
	.ZN(n424));
   AOI22_X1 U516 (.A1(n393),
	.A2(currIMM[15]),
	.B1(FE_OFN23_n394),
	.B2(MEM_DATA[15]),
	.ZN(n422));
   AOI22_X1 U517 (.A1(n393),
	.A2(currIMM[14]),
	.B1(FE_OFN23_n394),
	.B2(MEM_DATA[14]),
	.ZN(n423));
   AOI22_X1 U518 (.A1(FE_OFN19_n393),
	.A2(currIMM[10]),
	.B1(FE_OFN26_n394),
	.B2(MEM_DATA[10]),
	.ZN(n427));
   AOI22_X1 U519 (.A1(FE_OFN19_n393),
	.A2(currIMM[12]),
	.B1(FE_OFN25_n394),
	.B2(MEM_DATA[12]),
	.ZN(n425));
   AOI22_X1 U520 (.A1(n393),
	.A2(currIMM[11]),
	.B1(FE_OFN23_n394),
	.B2(MEM_DATA[11]),
	.ZN(n426));
   AOI22_X1 U521 (.A1(FE_OFN22_n393),
	.A2(currIMM[27]),
	.B1(FE_OFN28_n394),
	.B2(MEM_DATA[27]),
	.ZN(n409));
   AOI22_X1 U522 (.A1(FE_OFN22_n393),
	.A2(currIMM[26]),
	.B1(FE_OFN28_n394),
	.B2(MEM_DATA[26]),
	.ZN(n410));
   AOI22_X1 U523 (.A1(FE_OFN22_n393),
	.A2(currIMM[25]),
	.B1(FE_OFN28_n394),
	.B2(MEM_DATA[25]),
	.ZN(n411));
   AOI22_X1 U524 (.A1(FE_OFN22_n393),
	.A2(currIMM[24]),
	.B1(FE_OFN28_n394),
	.B2(MEM_DATA[24]),
	.ZN(n412));
   AOI22_X1 U525 (.A1(FE_OFN19_n393),
	.A2(currIMM[9]),
	.B1(FE_OFN23_n394),
	.B2(MEM_DATA[9]),
	.ZN(n392));
   AOI22_X1 U526 (.A1(FE_OFN22_n393),
	.A2(currIMM[23]),
	.B1(FE_OFN28_n394),
	.B2(MEM_DATA[23]),
	.ZN(n413));
   AOI22_X1 U527 (.A1(FE_OFN22_n393),
	.A2(currIMM[22]),
	.B1(FE_OFN28_n394),
	.B2(MEM_DATA[22]),
	.ZN(n414));
   AOI22_X1 U528 (.A1(FE_OFN22_n393),
	.A2(currIMM[21]),
	.B1(FE_OFN28_n394),
	.B2(MEM_DATA[21]),
	.ZN(n415));
   AOI22_X1 U529 (.A1(FE_OFN22_n393),
	.A2(currIMM[20]),
	.B1(FE_OFN28_n394),
	.B2(MEM_DATA[20]),
	.ZN(n416));
   AOI22_X1 U530 (.A1(FE_OFN20_n393),
	.A2(currIMM[1]),
	.B1(FE_OFN28_n394),
	.B2(MEM_DATA[1]),
	.ZN(n417));
   AOI22_X1 U531 (.A1(FE_OFN22_n393),
	.A2(currIMM[19]),
	.B1(FE_OFN28_n394),
	.B2(MEM_DATA[19]),
	.ZN(n418));
   AOI22_X1 U532 (.A1(FE_OFN19_n393),
	.A2(currIMM[16]),
	.B1(FE_OFN24_n394),
	.B2(MEM_DATA[16]),
	.ZN(n421));
   AOI22_X1 U533 (.A1(FE_OFN22_n393),
	.A2(currIMM[18]),
	.B1(FE_OFN28_n394),
	.B2(MEM_DATA[18]),
	.ZN(n419));
   AOI22_X1 U534 (.A1(FE_OFN39_ALU_OPA_SEL_c_2),
	.A2(MEM_WB_IN[19]),
	.B1(FE_OFN91_n432),
	.B2(currPC[19]),
	.ZN(n453));
   AOI22_X1 U535 (.A1(FE_OFN39_ALU_OPA_SEL_c_2),
	.A2(MEM_WB_IN[18]),
	.B1(FE_OFN91_n432),
	.B2(currPC[18]),
	.ZN(n454));
   AOI22_X1 U536 (.A1(FE_OFN39_ALU_OPA_SEL_c_2),
	.A2(MEM_WB_IN[17]),
	.B1(FE_OFN90_n432),
	.B2(currPC[17]),
	.ZN(n455));
   AOI22_X1 U537 (.A1(ALU_OPA_SEL[2]),
	.A2(MEM_WB_IN[16]),
	.B1(FE_OFN90_n432),
	.B2(currPC[16]),
	.ZN(n456));
   AOI22_X1 U538 (.A1(ALU_OPA_SEL[2]),
	.A2(MEM_WB_IN[15]),
	.B1(FE_OFN90_n432),
	.B2(currPC[15]),
	.ZN(n457));
   AOI22_X1 U539 (.A1(ALU_OPA_SEL[2]),
	.A2(MEM_WB_IN[14]),
	.B1(FE_OFN90_n432),
	.B2(currPC[14]),
	.ZN(n458));
   AOI22_X1 U540 (.A1(ALU_OPA_SEL[2]),
	.A2(MEM_WB_IN[13]),
	.B1(FE_OFN90_n432),
	.B2(currPC[13]),
	.ZN(n459));
   AOI22_X1 U541 (.A1(ALU_OPA_SEL[2]),
	.A2(MEM_WB_IN[12]),
	.B1(FE_OFN90_n432),
	.B2(currPC[12]),
	.ZN(n460));
   AOI22_X1 U542 (.A1(ALU_OPA_SEL[2]),
	.A2(MEM_WB_IN[11]),
	.B1(FE_OFN90_n432),
	.B2(currPC[11]),
	.ZN(n461));
   AOI22_X1 U543 (.A1(ALU_OPA_SEL[2]),
	.A2(MEM_WB_IN[10]),
	.B1(FE_OFN90_n432),
	.B2(currPC[10]),
	.ZN(n462));
   AOI22_X1 U544 (.A1(FE_OFN39_ALU_OPA_SEL_c_2),
	.A2(MEM_WB_IN[1]),
	.B1(FE_OFN90_n432),
	.B2(currPC[1]),
	.ZN(n452));
   OAI221_X1 U545 (.A(n463),
	.B1(n74),
	.B2(n429),
	.C1(n236),
	.C2(n430),
	.ZN(ALU_OPA[0]));
   AOI22_X1 U546 (.A1(ALU_OPA_SEL[2]),
	.A2(MEM_WB_IN[0]),
	.B1(n55),
	.B2(currPC[0]),
	.ZN(n463));
   NOR3_X1 U547 (.A1(ALU_OPA_SEL[1]),
	.A2(ALU_OPA_SEL[0]),
	.A3(ALU_OPA_SEL[2]),
	.ZN(n432));
   NOR3_X1 U548 (.A1(ALU_OPB_SEL[1]),
	.A2(ALU_OPB_SEL[2]),
	.A3(ALU_OPB_SEL[0]),
	.ZN(n394));
   AOI22_X1 U549 (.A1(FE_OFN22_n393),
	.A2(currIMM[30]),
	.B1(FE_OFN28_n394),
	.B2(MEM_DATA[30]),
	.ZN(n402));
   AOI22_X1 U550 (.A1(FE_OFN22_n393),
	.A2(currIMM[31]),
	.B1(FE_OFN28_n394),
	.B2(MEM_DATA[31]),
	.ZN(n401));
   AOI22_X1 U551 (.A1(FE_OFN22_n393),
	.A2(currIMM[29]),
	.B1(FE_OFN28_n394),
	.B2(MEM_DATA[29]),
	.ZN(n407));
   AOI22_X1 U552 (.A1(FE_OFN22_n393),
	.A2(currIMM[28]),
	.B1(FE_OFN28_n394),
	.B2(MEM_DATA[28]),
	.ZN(n408));
   AOI22_X1 U553 (.A1(FE_OFN19_n393),
	.A2(currIMM[8]),
	.B1(FE_OFN23_n394),
	.B2(MEM_DATA[8]),
	.ZN(n395));
   AOI22_X1 U554 (.A1(FE_OFN19_n393),
	.A2(currIMM[7]),
	.B1(FE_OFN23_n394),
	.B2(MEM_DATA[7]),
	.ZN(n396));
   AOI22_X1 U555 (.A1(FE_OFN20_n393),
	.A2(currIMM[6]),
	.B1(FE_OFN23_n394),
	.B2(MEM_DATA[6]),
	.ZN(n397));
   AOI22_X1 U556 (.A1(FE_OFN19_n393),
	.A2(currIMM[5]),
	.B1(FE_OFN23_n394),
	.B2(MEM_DATA[5]),
	.ZN(n398));
   AOI22_X1 U557 (.A1(n393),
	.A2(currIMM[4]),
	.B1(FE_OFN23_n394),
	.B2(MEM_DATA[4]),
	.ZN(n399));
   AOI22_X1 U558 (.A1(FE_OFN20_n393),
	.A2(currIMM[3]),
	.B1(FE_OFN27_n394),
	.B2(MEM_DATA[3]),
	.ZN(n400));
   AOI22_X1 U559 (.A1(FE_OFN19_n393),
	.A2(currIMM[0]),
	.B1(FE_OFN23_n394),
	.B2(MEM_DATA[0]),
	.ZN(n428));
   OAI221_X1 U560 (.A(n428),
	.B1(FE_DBTN0_n37),
	.B2(n236),
	.C1(n391),
	.C2(n204),
	.ZN(ALU_OPB[0]));
   INV_X1 U561 (.A(ALU_OPB_SEL[0]),
	.ZN(n172));
endmodule

module mem_unit (
	clk, 
	rst, 
	en, 
	ALU_OUT_IN, 
	MEM_DATA, 
	DRAM_OUT_IN, 
	DRAM_WR_IN, 
	DRAM_RD_IN, 
	RD_IN, 
	RD_OUT, 
	DRAM_WR, 
	DRAM_RD, 
	ALU_OUT, 
	DRAM_OUT, 
	DRAM_IN);
   input clk;
   input rst;
   input en;
   input [31:0] ALU_OUT_IN;
   input [31:0] MEM_DATA;
   input [31:0] DRAM_OUT_IN;
   input DRAM_WR_IN;
   input DRAM_RD_IN;
   input [4:0] RD_IN;
   output [4:0] RD_OUT;
   output DRAM_WR;
   output DRAM_RD;
   output [31:0] ALU_OUT;
   output [31:0] DRAM_OUT;
   output [31:0] DRAM_IN;

   // Internal wires
   wire FE_OFN58_n71;
   wire FE_OFN17_n72;
   wire n70;
   wire n71;
   wire n72;
   wire n73;
   wire n74;
   wire n75;
   wire n76;
   wire n77;
   wire n78;
   wire n79;
   wire n80;
   wire n81;
   wire n82;
   wire n83;
   wire n84;
   wire n85;
   wire n86;
   wire n87;
   wire n88;
   wire n89;
   wire n90;
   wire n91;
   wire n92;
   wire n93;
   wire n94;
   wire n95;
   wire n96;
   wire n97;
   wire n98;
   wire n99;
   wire n100;
   wire n101;
   wire n102;
   wire n103;
   wire n104;
   wire n105;
   wire n106;
   wire n107;
   wire n108;
   wire n109;
   wire n110;
   wire n111;
   wire n112;
   wire n113;
   wire n114;
   wire n115;
   wire n116;
   wire n117;
   wire n118;
   wire n119;
   wire n120;
   wire n121;
   wire n122;
   wire n123;
   wire n124;
   wire n125;
   wire n126;
   wire n127;
   wire n128;
   wire n129;
   wire n130;
   wire n131;
   wire n132;
   wire n133;
   wire n134;
   wire n135;
   wire n136;
   wire n137;
   wire n138;
   wire n139;
   wire n140;
   wire n1;
   wire n2;
   wire n3;
   wire n4;
   wire n18;
   wire n19;
   wire n20;
   wire n21;
   wire n22;
   wire n23;
   wire n24;
   wire n25;
   wire n26;
   wire n27;
   wire n28;
   wire n29;
   wire n30;
   wire n31;
   wire n32;
   wire n33;
   wire n34;
   wire n35;
   wire n36;
   wire n37;
   wire n38;
   wire n39;
   wire n40;
   wire n41;
   wire n42;
   wire n43;
   wire n44;
   wire n45;
   wire n46;
   wire n47;
   wire n48;
   wire n49;
   wire n50;
   wire n51;
   wire n52;
   wire n53;
   wire n54;
   wire n55;
   wire n56;
   wire n57;
   wire n58;
   wire n59;
   wire n60;
   wire n61;
   wire n62;
   wire n63;
   wire n64;
   wire n65;
   wire n66;
   wire n67;
   wire n68;
   wire n69;
   wire n141;
   wire n142;
   wire n143;
   wire n144;
   wire n145;
   wire n146;
   wire n147;
   wire n148;
   wire n149;
   wire n150;
   wire n151;
   wire n152;
   wire n153;
   wire n154;
   wire n155;
   wire n156;
   wire n157;

   assign DRAM_WR = DRAM_WR_IN ;
   assign DRAM_RD = DRAM_RD_IN ;
   assign DRAM_OUT[31] = DRAM_OUT_IN[31] ;
   assign DRAM_OUT[30] = DRAM_OUT_IN[30] ;
   assign DRAM_OUT[29] = DRAM_OUT_IN[29] ;
   assign DRAM_OUT[28] = DRAM_OUT_IN[28] ;
   assign DRAM_OUT[27] = DRAM_OUT_IN[27] ;
   assign DRAM_OUT[26] = DRAM_OUT_IN[26] ;
   assign DRAM_OUT[25] = DRAM_OUT_IN[25] ;
   assign DRAM_OUT[24] = DRAM_OUT_IN[24] ;
   assign DRAM_OUT[23] = DRAM_OUT_IN[23] ;
   assign DRAM_OUT[22] = DRAM_OUT_IN[22] ;
   assign DRAM_OUT[21] = DRAM_OUT_IN[21] ;
   assign DRAM_OUT[20] = DRAM_OUT_IN[20] ;
   assign DRAM_OUT[19] = DRAM_OUT_IN[19] ;
   assign DRAM_OUT[18] = DRAM_OUT_IN[18] ;
   assign DRAM_OUT[17] = DRAM_OUT_IN[17] ;
   assign DRAM_OUT[16] = DRAM_OUT_IN[16] ;
   assign DRAM_OUT[15] = DRAM_OUT_IN[15] ;
   assign DRAM_OUT[14] = DRAM_OUT_IN[14] ;
   assign DRAM_OUT[13] = DRAM_OUT_IN[13] ;
   assign DRAM_OUT[12] = DRAM_OUT_IN[12] ;
   assign DRAM_OUT[11] = DRAM_OUT_IN[11] ;
   assign DRAM_OUT[10] = DRAM_OUT_IN[10] ;
   assign DRAM_OUT[9] = DRAM_OUT_IN[9] ;
   assign DRAM_OUT[8] = DRAM_OUT_IN[8] ;
   assign DRAM_OUT[7] = DRAM_OUT_IN[7] ;
   assign DRAM_OUT[6] = DRAM_OUT_IN[6] ;
   assign DRAM_OUT[5] = DRAM_OUT_IN[5] ;
   assign DRAM_OUT[4] = DRAM_OUT_IN[4] ;
   assign DRAM_OUT[3] = DRAM_OUT_IN[3] ;
   assign DRAM_OUT[2] = DRAM_OUT_IN[2] ;
   assign DRAM_OUT[1] = DRAM_OUT_IN[1] ;
   assign DRAM_OUT[0] = DRAM_OUT_IN[0] ;

   CLKBUF_X3 FE_OFC58_n71 (.A(n71),
	.Z(FE_OFN58_n71));
   CLKBUF_X3 FE_OFC17_n72 (.A(n72),
	.Z(FE_OFN17_n72));
   DFF_X1 currALU_reg_29_ (.D(n19),
	.CK(clk),
	.Q(ALU_OUT[29]));
   DFF_X1 currALU_reg_28_ (.D(n20),
	.CK(clk),
	.Q(ALU_OUT[28]));
   DFF_X1 currALU_reg_27_ (.D(n21),
	.CK(clk),
	.Q(ALU_OUT[27]));
   DFF_X1 currALU_reg_26_ (.D(n22),
	.CK(clk),
	.Q(ALU_OUT[26]));
   DFF_X1 currALU_reg_25_ (.D(n23),
	.CK(clk),
	.Q(ALU_OUT[25]));
   DFF_X1 currALU_reg_24_ (.D(n24),
	.CK(clk),
	.Q(ALU_OUT[24]));
   DFF_X1 currALU_reg_23_ (.D(n25),
	.CK(clk),
	.Q(ALU_OUT[23]));
   DFF_X1 currALU_reg_22_ (.D(n26),
	.CK(clk),
	.Q(ALU_OUT[22]));
   DFF_X1 currALU_reg_21_ (.D(n27),
	.CK(clk),
	.Q(ALU_OUT[21]));
   DFF_X1 currALU_reg_20_ (.D(n28),
	.CK(clk),
	.Q(ALU_OUT[20]));
   DFF_X1 currALU_reg_19_ (.D(n29),
	.CK(clk),
	.Q(ALU_OUT[19]));
   DFF_X1 currALU_reg_18_ (.D(n30),
	.CK(clk),
	.Q(ALU_OUT[18]));
   DFF_X1 currALU_reg_17_ (.D(n31),
	.CK(clk),
	.Q(ALU_OUT[17]));
   DFF_X1 currALU_reg_16_ (.D(n32),
	.CK(clk),
	.Q(ALU_OUT[16]));
   DFF_X1 currALU_reg_15_ (.D(n33),
	.CK(clk),
	.Q(ALU_OUT[15]));
   DFF_X1 currALU_reg_14_ (.D(n34),
	.CK(clk),
	.Q(ALU_OUT[14]));
   DFF_X1 currALU_reg_13_ (.D(n35),
	.CK(clk),
	.Q(ALU_OUT[13]));
   DFF_X1 currALU_reg_12_ (.D(n36),
	.CK(clk),
	.Q(ALU_OUT[12]));
   DFF_X1 currALU_reg_11_ (.D(n37),
	.CK(clk),
	.Q(ALU_OUT[11]));
   DFF_X1 currALU_reg_10_ (.D(n38),
	.CK(clk),
	.Q(ALU_OUT[10]));
   DFF_X1 currALU_reg_9_ (.D(n39),
	.CK(clk),
	.Q(ALU_OUT[9]));
   DFF_X1 currALU_reg_8_ (.D(n40),
	.CK(clk),
	.Q(ALU_OUT[8]));
   DFF_X1 currALU_reg_7_ (.D(n41),
	.CK(clk),
	.Q(ALU_OUT[7]));
   DFF_X1 currALU_reg_6_ (.D(n42),
	.CK(clk),
	.Q(ALU_OUT[6]));
   DFF_X1 currALU_reg_5_ (.D(n43),
	.CK(clk),
	.Q(ALU_OUT[5]));
   DFF_X1 currALU_reg_4_ (.D(n44),
	.CK(clk),
	.Q(ALU_OUT[4]));
   DFF_X1 currALU_reg_3_ (.D(n45),
	.CK(clk),
	.Q(ALU_OUT[3]));
   DFF_X1 currALU_reg_2_ (.D(n46),
	.CK(clk),
	.Q(ALU_OUT[2]));
   DFF_X1 currALU_reg_1_ (.D(n47),
	.CK(clk),
	.Q(ALU_OUT[1]));
   DFF_X1 currALU_reg_0_ (.D(n48),
	.CK(clk),
	.Q(ALU_OUT[0]));
   DFF_X1 currMEM_DATA_reg_31_ (.D(n55),
	.CK(clk),
	.Q(DRAM_IN[31]));
   DFF_X1 currMEM_DATA_reg_30_ (.D(n56),
	.CK(clk),
	.Q(DRAM_IN[30]));
   DFF_X1 currMEM_DATA_reg_29_ (.D(n57),
	.CK(clk),
	.Q(DRAM_IN[29]));
   DFF_X1 currMEM_DATA_reg_28_ (.D(n58),
	.CK(clk),
	.Q(DRAM_IN[28]));
   DFF_X1 currMEM_DATA_reg_27_ (.D(n59),
	.CK(clk),
	.Q(DRAM_IN[27]));
   DFF_X1 currMEM_DATA_reg_26_ (.D(n60),
	.CK(clk),
	.Q(DRAM_IN[26]));
   DFF_X1 currMEM_DATA_reg_25_ (.D(n61),
	.CK(clk),
	.Q(DRAM_IN[25]));
   DFF_X1 currMEM_DATA_reg_24_ (.D(n62),
	.CK(clk),
	.Q(DRAM_IN[24]));
   DFF_X1 currMEM_DATA_reg_23_ (.D(n63),
	.CK(clk),
	.Q(DRAM_IN[23]));
   DFF_X1 currMEM_DATA_reg_22_ (.D(n64),
	.CK(clk),
	.Q(DRAM_IN[22]));
   DFF_X1 currMEM_DATA_reg_21_ (.D(n65),
	.CK(clk),
	.Q(DRAM_IN[21]));
   DFF_X1 currMEM_DATA_reg_20_ (.D(n66),
	.CK(clk),
	.Q(DRAM_IN[20]));
   DFF_X1 currMEM_DATA_reg_19_ (.D(n67),
	.CK(clk),
	.Q(DRAM_IN[19]));
   DFF_X1 currMEM_DATA_reg_18_ (.D(n68),
	.CK(clk),
	.Q(DRAM_IN[18]));
   DFF_X1 currMEM_DATA_reg_17_ (.D(n69),
	.CK(clk),
	.Q(DRAM_IN[17]));
   DFF_X1 currMEM_DATA_reg_16_ (.D(n141),
	.CK(clk),
	.Q(DRAM_IN[16]));
   DFF_X1 currMEM_DATA_reg_15_ (.D(n142),
	.CK(clk),
	.Q(DRAM_IN[15]));
   DFF_X1 currMEM_DATA_reg_14_ (.D(n143),
	.CK(clk),
	.Q(DRAM_IN[14]));
   DFF_X1 currMEM_DATA_reg_13_ (.D(n144),
	.CK(clk),
	.Q(DRAM_IN[13]));
   DFF_X1 currMEM_DATA_reg_12_ (.D(n145),
	.CK(clk),
	.Q(DRAM_IN[12]));
   DFF_X1 currMEM_DATA_reg_11_ (.D(n146),
	.CK(clk),
	.Q(DRAM_IN[11]));
   DFF_X1 currMEM_DATA_reg_10_ (.D(n147),
	.CK(clk),
	.Q(DRAM_IN[10]));
   DFF_X1 currMEM_DATA_reg_9_ (.D(n148),
	.CK(clk),
	.Q(DRAM_IN[9]));
   DFF_X1 currMEM_DATA_reg_8_ (.D(n149),
	.CK(clk),
	.Q(DRAM_IN[8]));
   DFF_X1 currMEM_DATA_reg_7_ (.D(n150),
	.CK(clk),
	.Q(DRAM_IN[7]));
   DFF_X1 currMEM_DATA_reg_6_ (.D(n151),
	.CK(clk),
	.Q(DRAM_IN[6]));
   DFF_X1 currMEM_DATA_reg_5_ (.D(n152),
	.CK(clk),
	.Q(DRAM_IN[5]));
   DFF_X1 currMEM_DATA_reg_4_ (.D(n153),
	.CK(clk),
	.Q(DRAM_IN[4]));
   DFF_X1 currMEM_DATA_reg_3_ (.D(n154),
	.CK(clk),
	.Q(DRAM_IN[3]));
   DFF_X1 currMEM_DATA_reg_2_ (.D(n155),
	.CK(clk),
	.Q(DRAM_IN[2]));
   DFF_X1 currMEM_DATA_reg_1_ (.D(n156),
	.CK(clk),
	.Q(DRAM_IN[1]));
   DFF_X1 currMEM_DATA_reg_0_ (.D(n157),
	.CK(clk),
	.Q(DRAM_IN[0]));
   DFF_X1 currALU_reg_30_ (.D(n18),
	.CK(clk),
	.Q(ALU_OUT[30]));
   DFF_X1 currALU_reg_31_ (.D(n49),
	.CK(clk),
	.Q(ALU_OUT[31]));
   DFF_X1 currRD_reg_1_ (.D(n53),
	.CK(clk),
	.Q(RD_OUT[1]));
   DFF_X1 currRD_reg_0_ (.D(n54),
	.CK(clk),
	.Q(RD_OUT[0]));
   DFF_X1 currRD_reg_2_ (.D(n52),
	.CK(clk),
	.Q(RD_OUT[2]),
	.QN(n3));
   DFF_X1 currRD_reg_4_ (.D(n50),
	.CK(clk),
	.Q(RD_OUT[4]),
	.QN(n1));
   DFF_X1 currRD_reg_3_ (.D(n51),
	.CK(clk),
	.Q(RD_OUT[3]));
   INV_X1 U3 (.A(n1),
	.ZN(n2));
   INV_X1 U4 (.A(n3),
	.ZN(n4));
   INV_X1 U17 (.A(n134),
	.ZN(n18));
   AOI22_X1 U18 (.A1(ALU_OUT_IN[30]),
	.A2(FE_OFN58_n71),
	.B1(ALU_OUT[30]),
	.B2(FE_OFN17_n72),
	.ZN(n134));
   INV_X1 U19 (.A(n133),
	.ZN(n19));
   AOI22_X1 U20 (.A1(ALU_OUT_IN[29]),
	.A2(FE_OFN58_n71),
	.B1(ALU_OUT[29]),
	.B2(FE_OFN17_n72),
	.ZN(n133));
   INV_X1 U21 (.A(n132),
	.ZN(n20));
   AOI22_X1 U22 (.A1(ALU_OUT_IN[28]),
	.A2(FE_OFN58_n71),
	.B1(ALU_OUT[28]),
	.B2(FE_OFN17_n72),
	.ZN(n132));
   INV_X1 U23 (.A(n131),
	.ZN(n21));
   AOI22_X1 U24 (.A1(ALU_OUT_IN[27]),
	.A2(FE_OFN58_n71),
	.B1(ALU_OUT[27]),
	.B2(FE_OFN17_n72),
	.ZN(n131));
   INV_X1 U25 (.A(n130),
	.ZN(n22));
   AOI22_X1 U26 (.A1(ALU_OUT_IN[26]),
	.A2(FE_OFN58_n71),
	.B1(ALU_OUT[26]),
	.B2(FE_OFN17_n72),
	.ZN(n130));
   INV_X1 U27 (.A(n124),
	.ZN(n28));
   AOI22_X1 U28 (.A1(ALU_OUT_IN[20]),
	.A2(FE_OFN58_n71),
	.B1(ALU_OUT[20]),
	.B2(FE_OFN17_n72),
	.ZN(n124));
   INV_X1 U29 (.A(n125),
	.ZN(n27));
   AOI22_X1 U30 (.A1(ALU_OUT_IN[21]),
	.A2(FE_OFN58_n71),
	.B1(ALU_OUT[21]),
	.B2(FE_OFN17_n72),
	.ZN(n125));
   INV_X1 U31 (.A(n126),
	.ZN(n26));
   AOI22_X1 U32 (.A1(ALU_OUT_IN[22]),
	.A2(FE_OFN58_n71),
	.B1(ALU_OUT[22]),
	.B2(FE_OFN17_n72),
	.ZN(n126));
   INV_X1 U33 (.A(n129),
	.ZN(n23));
   AOI22_X1 U34 (.A1(ALU_OUT_IN[25]),
	.A2(FE_OFN58_n71),
	.B1(ALU_OUT[25]),
	.B2(FE_OFN17_n72),
	.ZN(n129));
   INV_X1 U35 (.A(n128),
	.ZN(n24));
   AOI22_X1 U36 (.A1(ALU_OUT_IN[24]),
	.A2(FE_OFN58_n71),
	.B1(ALU_OUT[24]),
	.B2(FE_OFN17_n72),
	.ZN(n128));
   INV_X1 U37 (.A(n127),
	.ZN(n25));
   AOI22_X1 U38 (.A1(ALU_OUT_IN[23]),
	.A2(FE_OFN58_n71),
	.B1(ALU_OUT[23]),
	.B2(FE_OFN17_n72),
	.ZN(n127));
   INV_X1 U39 (.A(n116),
	.ZN(n36));
   AOI22_X1 U40 (.A1(ALU_OUT_IN[12]),
	.A2(FE_OFN58_n71),
	.B1(ALU_OUT[12]),
	.B2(FE_OFN17_n72),
	.ZN(n116));
   INV_X1 U41 (.A(n117),
	.ZN(n35));
   AOI22_X1 U42 (.A1(ALU_OUT_IN[13]),
	.A2(FE_OFN58_n71),
	.B1(ALU_OUT[13]),
	.B2(FE_OFN17_n72),
	.ZN(n117));
   INV_X1 U43 (.A(n118),
	.ZN(n34));
   AOI22_X1 U44 (.A1(ALU_OUT_IN[14]),
	.A2(FE_OFN58_n71),
	.B1(ALU_OUT[14]),
	.B2(FE_OFN17_n72),
	.ZN(n118));
   INV_X1 U45 (.A(n119),
	.ZN(n33));
   AOI22_X1 U46 (.A1(ALU_OUT_IN[15]),
	.A2(FE_OFN58_n71),
	.B1(ALU_OUT[15]),
	.B2(FE_OFN17_n72),
	.ZN(n119));
   INV_X1 U47 (.A(n120),
	.ZN(n32));
   AOI22_X1 U48 (.A1(ALU_OUT_IN[16]),
	.A2(FE_OFN58_n71),
	.B1(ALU_OUT[16]),
	.B2(FE_OFN17_n72),
	.ZN(n120));
   INV_X1 U49 (.A(n121),
	.ZN(n31));
   AOI22_X1 U50 (.A1(ALU_OUT_IN[17]),
	.A2(FE_OFN58_n71),
	.B1(ALU_OUT[17]),
	.B2(FE_OFN17_n72),
	.ZN(n121));
   INV_X1 U51 (.A(n122),
	.ZN(n30));
   AOI22_X1 U52 (.A1(ALU_OUT_IN[18]),
	.A2(FE_OFN58_n71),
	.B1(ALU_OUT[18]),
	.B2(FE_OFN17_n72),
	.ZN(n122));
   INV_X1 U53 (.A(n123),
	.ZN(n29));
   AOI22_X1 U54 (.A1(ALU_OUT_IN[19]),
	.A2(FE_OFN58_n71),
	.B1(ALU_OUT[19]),
	.B2(FE_OFN17_n72),
	.ZN(n123));
   INV_X1 U55 (.A(n104),
	.ZN(n48));
   AOI22_X1 U56 (.A1(ALU_OUT_IN[0]),
	.A2(FE_OFN58_n71),
	.B1(ALU_OUT[0]),
	.B2(FE_OFN17_n72),
	.ZN(n104));
   INV_X1 U57 (.A(n106),
	.ZN(n46));
   AOI22_X1 U58 (.A1(ALU_OUT_IN[2]),
	.A2(FE_OFN58_n71),
	.B1(ALU_OUT[2]),
	.B2(FE_OFN17_n72),
	.ZN(n106));
   INV_X1 U59 (.A(n107),
	.ZN(n45));
   AOI22_X1 U60 (.A1(ALU_OUT_IN[3]),
	.A2(FE_OFN58_n71),
	.B1(ALU_OUT[3]),
	.B2(FE_OFN17_n72),
	.ZN(n107));
   INV_X1 U61 (.A(n108),
	.ZN(n44));
   AOI22_X1 U62 (.A1(ALU_OUT_IN[4]),
	.A2(FE_OFN58_n71),
	.B1(ALU_OUT[4]),
	.B2(FE_OFN17_n72),
	.ZN(n108));
   INV_X1 U63 (.A(n109),
	.ZN(n43));
   AOI22_X1 U64 (.A1(ALU_OUT_IN[5]),
	.A2(FE_OFN58_n71),
	.B1(ALU_OUT[5]),
	.B2(FE_OFN17_n72),
	.ZN(n109));
   INV_X1 U65 (.A(n110),
	.ZN(n42));
   AOI22_X1 U66 (.A1(ALU_OUT_IN[6]),
	.A2(FE_OFN58_n71),
	.B1(ALU_OUT[6]),
	.B2(FE_OFN17_n72),
	.ZN(n110));
   INV_X1 U67 (.A(n111),
	.ZN(n41));
   AOI22_X1 U68 (.A1(ALU_OUT_IN[7]),
	.A2(FE_OFN58_n71),
	.B1(ALU_OUT[7]),
	.B2(FE_OFN17_n72),
	.ZN(n111));
   INV_X1 U69 (.A(n114),
	.ZN(n38));
   AOI22_X1 U70 (.A1(ALU_OUT_IN[10]),
	.A2(FE_OFN58_n71),
	.B1(ALU_OUT[10]),
	.B2(FE_OFN17_n72),
	.ZN(n114));
   INV_X1 U71 (.A(n105),
	.ZN(n47));
   AOI22_X1 U72 (.A1(ALU_OUT_IN[1]),
	.A2(FE_OFN58_n71),
	.B1(ALU_OUT[1]),
	.B2(FE_OFN17_n72),
	.ZN(n105));
   INV_X1 U73 (.A(n112),
	.ZN(n40));
   AOI22_X1 U74 (.A1(ALU_OUT_IN[8]),
	.A2(FE_OFN58_n71),
	.B1(ALU_OUT[8]),
	.B2(FE_OFN17_n72),
	.ZN(n112));
   INV_X1 U75 (.A(n113),
	.ZN(n39));
   AOI22_X1 U76 (.A1(ALU_OUT_IN[9]),
	.A2(FE_OFN58_n71),
	.B1(ALU_OUT[9]),
	.B2(FE_OFN17_n72),
	.ZN(n113));
   INV_X1 U77 (.A(n115),
	.ZN(n37));
   AOI22_X1 U78 (.A1(ALU_OUT_IN[11]),
	.A2(FE_OFN58_n71),
	.B1(ALU_OUT[11]),
	.B2(FE_OFN17_n72),
	.ZN(n115));
   NOR2_X1 U79 (.A1(en),
	.A2(rst),
	.ZN(n72));
   NOR2_X1 U81 (.A1(n72),
	.A2(rst),
	.ZN(n71));
   INV_X1 U82 (.A(n139),
	.ZN(n51));
   AOI22_X1 U83 (.A1(RD_IN[3]),
	.A2(n71),
	.B1(RD_OUT[3]),
	.B2(n72),
	.ZN(n139));
   INV_X1 U84 (.A(n140),
	.ZN(n50));
   AOI22_X1 U85 (.A1(RD_IN[4]),
	.A2(n71),
	.B1(n2),
	.B2(n72),
	.ZN(n140));
   INV_X1 U86 (.A(n136),
	.ZN(n54));
   INV_X1 U87 (.A(n137),
	.ZN(n53));
   INV_X1 U88 (.A(n70),
	.ZN(n157));
   AOI22_X1 U89 (.A1(MEM_DATA[0]),
	.A2(FE_OFN58_n71),
	.B1(DRAM_IN[0]),
	.B2(FE_OFN17_n72),
	.ZN(n70));
   INV_X1 U90 (.A(n73),
	.ZN(n156));
   AOI22_X1 U91 (.A1(MEM_DATA[1]),
	.A2(FE_OFN58_n71),
	.B1(DRAM_IN[1]),
	.B2(FE_OFN17_n72),
	.ZN(n73));
   INV_X1 U92 (.A(n74),
	.ZN(n155));
   AOI22_X1 U93 (.A1(MEM_DATA[2]),
	.A2(FE_OFN58_n71),
	.B1(DRAM_IN[2]),
	.B2(FE_OFN17_n72),
	.ZN(n74));
   INV_X1 U94 (.A(n75),
	.ZN(n154));
   AOI22_X1 U95 (.A1(MEM_DATA[3]),
	.A2(FE_OFN58_n71),
	.B1(DRAM_IN[3]),
	.B2(FE_OFN17_n72),
	.ZN(n75));
   INV_X1 U96 (.A(n76),
	.ZN(n153));
   AOI22_X1 U97 (.A1(MEM_DATA[4]),
	.A2(FE_OFN58_n71),
	.B1(DRAM_IN[4]),
	.B2(FE_OFN17_n72),
	.ZN(n76));
   INV_X1 U98 (.A(n77),
	.ZN(n152));
   AOI22_X1 U99 (.A1(MEM_DATA[5]),
	.A2(FE_OFN58_n71),
	.B1(DRAM_IN[5]),
	.B2(FE_OFN17_n72),
	.ZN(n77));
   INV_X1 U100 (.A(n78),
	.ZN(n151));
   AOI22_X1 U101 (.A1(MEM_DATA[6]),
	.A2(FE_OFN58_n71),
	.B1(DRAM_IN[6]),
	.B2(FE_OFN17_n72),
	.ZN(n78));
   INV_X1 U102 (.A(n79),
	.ZN(n150));
   AOI22_X1 U103 (.A1(MEM_DATA[7]),
	.A2(FE_OFN58_n71),
	.B1(DRAM_IN[7]),
	.B2(FE_OFN17_n72),
	.ZN(n79));
   INV_X1 U104 (.A(n80),
	.ZN(n149));
   AOI22_X1 U105 (.A1(MEM_DATA[8]),
	.A2(FE_OFN58_n71),
	.B1(DRAM_IN[8]),
	.B2(FE_OFN17_n72),
	.ZN(n80));
   INV_X1 U106 (.A(n81),
	.ZN(n148));
   AOI22_X1 U107 (.A1(MEM_DATA[9]),
	.A2(FE_OFN58_n71),
	.B1(DRAM_IN[9]),
	.B2(FE_OFN17_n72),
	.ZN(n81));
   INV_X1 U108 (.A(n82),
	.ZN(n147));
   AOI22_X1 U109 (.A1(MEM_DATA[10]),
	.A2(FE_OFN58_n71),
	.B1(DRAM_IN[10]),
	.B2(FE_OFN17_n72),
	.ZN(n82));
   INV_X1 U110 (.A(n83),
	.ZN(n146));
   AOI22_X1 U111 (.A1(MEM_DATA[11]),
	.A2(n71),
	.B1(DRAM_IN[11]),
	.B2(n72),
	.ZN(n83));
   INV_X1 U112 (.A(n84),
	.ZN(n145));
   AOI22_X1 U113 (.A1(MEM_DATA[12]),
	.A2(FE_OFN58_n71),
	.B1(DRAM_IN[12]),
	.B2(FE_OFN17_n72),
	.ZN(n84));
   INV_X1 U114 (.A(n85),
	.ZN(n144));
   AOI22_X1 U115 (.A1(MEM_DATA[13]),
	.A2(FE_OFN58_n71),
	.B1(DRAM_IN[13]),
	.B2(FE_OFN17_n72),
	.ZN(n85));
   INV_X1 U116 (.A(n86),
	.ZN(n143));
   AOI22_X1 U117 (.A1(MEM_DATA[14]),
	.A2(n71),
	.B1(DRAM_IN[14]),
	.B2(FE_OFN17_n72),
	.ZN(n86));
   INV_X1 U118 (.A(n87),
	.ZN(n142));
   AOI22_X1 U119 (.A1(MEM_DATA[15]),
	.A2(FE_OFN58_n71),
	.B1(DRAM_IN[15]),
	.B2(FE_OFN17_n72),
	.ZN(n87));
   INV_X1 U120 (.A(n88),
	.ZN(n141));
   AOI22_X1 U121 (.A1(MEM_DATA[16]),
	.A2(FE_OFN58_n71),
	.B1(DRAM_IN[16]),
	.B2(FE_OFN17_n72),
	.ZN(n88));
   INV_X1 U122 (.A(n89),
	.ZN(n69));
   AOI22_X1 U123 (.A1(MEM_DATA[17]),
	.A2(FE_OFN58_n71),
	.B1(DRAM_IN[17]),
	.B2(FE_OFN17_n72),
	.ZN(n89));
   INV_X1 U124 (.A(n90),
	.ZN(n68));
   AOI22_X1 U125 (.A1(MEM_DATA[18]),
	.A2(FE_OFN58_n71),
	.B1(DRAM_IN[18]),
	.B2(FE_OFN17_n72),
	.ZN(n90));
   INV_X1 U126 (.A(n91),
	.ZN(n67));
   AOI22_X1 U127 (.A1(MEM_DATA[19]),
	.A2(FE_OFN58_n71),
	.B1(DRAM_IN[19]),
	.B2(FE_OFN17_n72),
	.ZN(n91));
   INV_X1 U128 (.A(n92),
	.ZN(n66));
   AOI22_X1 U129 (.A1(MEM_DATA[20]),
	.A2(FE_OFN58_n71),
	.B1(DRAM_IN[20]),
	.B2(FE_OFN17_n72),
	.ZN(n92));
   INV_X1 U130 (.A(n93),
	.ZN(n65));
   AOI22_X1 U131 (.A1(MEM_DATA[21]),
	.A2(FE_OFN58_n71),
	.B1(DRAM_IN[21]),
	.B2(FE_OFN17_n72),
	.ZN(n93));
   INV_X1 U132 (.A(n94),
	.ZN(n64));
   AOI22_X1 U133 (.A1(MEM_DATA[22]),
	.A2(FE_OFN58_n71),
	.B1(DRAM_IN[22]),
	.B2(FE_OFN17_n72),
	.ZN(n94));
   INV_X1 U134 (.A(n95),
	.ZN(n63));
   AOI22_X1 U135 (.A1(MEM_DATA[23]),
	.A2(FE_OFN58_n71),
	.B1(DRAM_IN[23]),
	.B2(FE_OFN17_n72),
	.ZN(n95));
   INV_X1 U136 (.A(n96),
	.ZN(n62));
   AOI22_X1 U137 (.A1(MEM_DATA[24]),
	.A2(FE_OFN58_n71),
	.B1(DRAM_IN[24]),
	.B2(FE_OFN17_n72),
	.ZN(n96));
   INV_X1 U138 (.A(n97),
	.ZN(n61));
   AOI22_X1 U139 (.A1(MEM_DATA[25]),
	.A2(FE_OFN58_n71),
	.B1(DRAM_IN[25]),
	.B2(FE_OFN17_n72),
	.ZN(n97));
   INV_X1 U140 (.A(n98),
	.ZN(n60));
   AOI22_X1 U141 (.A1(MEM_DATA[26]),
	.A2(FE_OFN58_n71),
	.B1(DRAM_IN[26]),
	.B2(FE_OFN17_n72),
	.ZN(n98));
   INV_X1 U142 (.A(n99),
	.ZN(n59));
   AOI22_X1 U143 (.A1(MEM_DATA[27]),
	.A2(FE_OFN58_n71),
	.B1(DRAM_IN[27]),
	.B2(FE_OFN17_n72),
	.ZN(n99));
   INV_X1 U144 (.A(n100),
	.ZN(n58));
   AOI22_X1 U145 (.A1(MEM_DATA[28]),
	.A2(FE_OFN58_n71),
	.B1(DRAM_IN[28]),
	.B2(FE_OFN17_n72),
	.ZN(n100));
   INV_X1 U146 (.A(n101),
	.ZN(n57));
   AOI22_X1 U147 (.A1(MEM_DATA[29]),
	.A2(FE_OFN58_n71),
	.B1(DRAM_IN[29]),
	.B2(FE_OFN17_n72),
	.ZN(n101));
   INV_X1 U148 (.A(n102),
	.ZN(n56));
   AOI22_X1 U149 (.A1(MEM_DATA[30]),
	.A2(FE_OFN58_n71),
	.B1(DRAM_IN[30]),
	.B2(FE_OFN17_n72),
	.ZN(n102));
   INV_X1 U150 (.A(n103),
	.ZN(n55));
   AOI22_X1 U151 (.A1(MEM_DATA[31]),
	.A2(FE_OFN58_n71),
	.B1(DRAM_IN[31]),
	.B2(FE_OFN17_n72),
	.ZN(n103));
   INV_X1 U152 (.A(n138),
	.ZN(n52));
   AOI22_X1 U153 (.A1(RD_IN[0]),
	.A2(n71),
	.B1(RD_OUT[0]),
	.B2(n72),
	.ZN(n136));
   AOI22_X1 U154 (.A1(RD_IN[2]),
	.A2(n71),
	.B1(n4),
	.B2(n72),
	.ZN(n138));
   AOI22_X1 U155 (.A1(RD_IN[1]),
	.A2(n71),
	.B1(RD_OUT[1]),
	.B2(n72),
	.ZN(n137));
   AOI22_X1 U156 (.A1(ALU_OUT_IN[31]),
	.A2(FE_OFN58_n71),
	.B1(ALU_OUT[31]),
	.B2(FE_OFN17_n72),
	.ZN(n135));
   INV_X1 U157 (.A(n135),
	.ZN(n49));
endmodule

module wb_unit (
	clk, 
	rst, 
	en, 
	RD_IN, 
	ALU_OUT, 
	DRAM_OUT, 
	MUX_SEL, 
	RD_OUT, 
	WB_OUT);
   input clk;
   input rst;
   input en;
   input [4:0] RD_IN;
   input [31:0] ALU_OUT;
   input [31:0] DRAM_OUT;
   input MUX_SEL;
   output [4:0] RD_OUT;
   output [31:0] WB_OUT;

   // Internal wires
   wire FE_OFN57_n105;
   wire FE_OFN41_MUX_SEL_WB_c;
   wire FE_OFN16_n104;
   wire FE_OFN15_n104;
   wire n103;
   wire n104;
   wire n105;
   wire n106;
   wire n107;
   wire n108;
   wire n109;
   wire n110;
   wire n111;
   wire n112;
   wire n113;
   wire n114;
   wire n115;
   wire n116;
   wire n117;
   wire n118;
   wire n119;
   wire n120;
   wire n121;
   wire n122;
   wire n123;
   wire n124;
   wire n125;
   wire n126;
   wire n127;
   wire n128;
   wire n129;
   wire n130;
   wire n131;
   wire n132;
   wire n133;
   wire n134;
   wire n135;
   wire n136;
   wire n137;
   wire n138;
   wire n139;
   wire n140;
   wire n141;
   wire n142;
   wire n143;
   wire n144;
   wire n145;
   wire n146;
   wire n147;
   wire n148;
   wire n149;
   wire n150;
   wire n151;
   wire n152;
   wire n153;
   wire n154;
   wire n155;
   wire n156;
   wire n157;
   wire n158;
   wire n159;
   wire n160;
   wire n161;
   wire n162;
   wire n163;
   wire n164;
   wire n165;
   wire n166;
   wire n167;
   wire n168;
   wire n169;
   wire n170;
   wire n171;
   wire n172;
   wire n173;
   wire n174;
   wire n175;
   wire n176;
   wire n177;
   wire n178;
   wire n179;
   wire n180;
   wire n181;
   wire n182;
   wire n183;
   wire n184;
   wire n185;
   wire n186;
   wire n187;
   wire n188;
   wire n189;
   wire n190;
   wire n191;
   wire n192;
   wire n193;
   wire n194;
   wire n195;
   wire n196;
   wire n197;
   wire n198;
   wire n199;
   wire n200;
   wire n201;
   wire n202;
   wire n203;
   wire n204;
   wire n205;
   wire n1;
   wire n2;
   wire n3;
   wire n4;
   wire n27;
   wire n28;
   wire n29;
   wire n30;
   wire n31;
   wire n32;
   wire n34;
   wire n36;
   wire n38;
   wire n40;
   wire n42;
   wire n44;
   wire n46;
   wire n48;
   wire n50;
   wire n52;
   wire n54;
   wire n56;
   wire n58;
   wire n60;
   wire n62;
   wire n64;
   wire n66;
   wire n68;
   wire n70;
   wire n72;
   wire n74;
   wire n76;
   wire n78;
   wire n80;
   wire n82;
   wire n84;
   wire n86;
   wire n88;
   wire n90;
   wire n92;
   wire n94;
   wire n96;
   wire n97;
   wire n98;
   wire n99;
   wire n100;
   wire n101;
   wire n102;
   wire n206;
   wire n207;
   wire n208;
   wire n209;
   wire n210;
   wire n211;
   wire n212;
   wire n213;
   wire n214;
   wire n215;
   wire n216;
   wire n217;
   wire n218;
   wire n219;
   wire n220;
   wire n221;
   wire n222;
   wire n223;
   wire n224;
   wire n225;
   wire n226;
   wire n227;
   wire n228;
   wire n229;
   wire n230;
   wire n231;
   wire [31:0] currALU;
   wire [31:0] currMEM;

   CLKBUF_X3 FE_OFC57_n105 (.A(n105),
	.Z(FE_OFN57_n105));
   BUF_X1 FE_OFC41_MUX_SEL_WB_c (.A(MUX_SEL),
	.Z(FE_OFN41_MUX_SEL_WB_c));
   BUF_X1 FE_OFC16_n104 (.A(FE_OFN15_n104),
	.Z(FE_OFN16_n104));
   BUF_X2 FE_OFC15_n104 (.A(n104),
	.Z(FE_OFN15_n104));
   DFF_X1 currALU_reg_31_ (.D(n34),
	.CK(clk),
	.Q(currALU[31]));
   DFF_X1 currALU_reg_30_ (.D(n36),
	.CK(clk),
	.Q(currALU[30]));
   DFF_X1 currALU_reg_29_ (.D(n38),
	.CK(clk),
	.Q(currALU[29]));
   DFF_X1 currALU_reg_28_ (.D(n40),
	.CK(clk),
	.Q(currALU[28]));
   DFF_X1 currALU_reg_27_ (.D(n42),
	.CK(clk),
	.Q(currALU[27]));
   DFF_X1 currALU_reg_26_ (.D(n44),
	.CK(clk),
	.Q(currALU[26]));
   DFF_X1 currALU_reg_25_ (.D(n46),
	.CK(clk),
	.Q(currALU[25]));
   DFF_X1 currALU_reg_24_ (.D(n48),
	.CK(clk),
	.Q(currALU[24]));
   DFF_X1 currALU_reg_23_ (.D(n50),
	.CK(clk),
	.Q(currALU[23]));
   DFF_X1 currALU_reg_22_ (.D(n52),
	.CK(clk),
	.Q(currALU[22]));
   DFF_X1 currALU_reg_21_ (.D(n54),
	.CK(clk),
	.Q(currALU[21]));
   DFF_X1 currALU_reg_20_ (.D(n56),
	.CK(clk),
	.Q(currALU[20]));
   DFF_X1 currALU_reg_19_ (.D(n58),
	.CK(clk),
	.Q(currALU[19]));
   DFF_X1 currALU_reg_18_ (.D(n60),
	.CK(clk),
	.Q(currALU[18]));
   DFF_X1 currALU_reg_17_ (.D(n62),
	.CK(clk),
	.Q(currALU[17]));
   DFF_X1 currALU_reg_16_ (.D(n64),
	.CK(clk),
	.Q(currALU[16]));
   DFF_X1 currALU_reg_15_ (.D(n66),
	.CK(clk),
	.Q(currALU[15]));
   DFF_X1 currALU_reg_14_ (.D(n68),
	.CK(clk),
	.Q(currALU[14]));
   DFF_X1 currALU_reg_13_ (.D(n70),
	.CK(clk),
	.Q(currALU[13]));
   DFF_X1 currALU_reg_12_ (.D(n72),
	.CK(clk),
	.Q(currALU[12]));
   DFF_X1 currALU_reg_11_ (.D(n74),
	.CK(clk),
	.Q(currALU[11]));
   DFF_X1 currALU_reg_10_ (.D(n76),
	.CK(clk),
	.Q(currALU[10]));
   DFF_X1 currALU_reg_9_ (.D(n78),
	.CK(clk),
	.Q(currALU[9]));
   DFF_X1 currALU_reg_8_ (.D(n80),
	.CK(clk),
	.Q(currALU[8]));
   DFF_X1 currALU_reg_7_ (.D(n82),
	.CK(clk),
	.Q(currALU[7]));
   DFF_X1 currALU_reg_6_ (.D(n84),
	.CK(clk),
	.Q(currALU[6]));
   DFF_X1 currALU_reg_5_ (.D(n86),
	.CK(clk),
	.Q(currALU[5]));
   DFF_X1 currALU_reg_4_ (.D(n88),
	.CK(clk),
	.Q(currALU[4]));
   DFF_X1 currALU_reg_3_ (.D(n90),
	.CK(clk),
	.Q(currALU[3]));
   DFF_X1 currALU_reg_2_ (.D(n92),
	.CK(clk),
	.Q(currALU[2]));
   DFF_X1 currALU_reg_1_ (.D(n94),
	.CK(clk),
	.Q(currALU[1]));
   DFF_X1 currALU_reg_0_ (.D(n96),
	.CK(clk),
	.Q(currALU[0]));
   DFF_X1 currMEM_reg_31_ (.D(n97),
	.CK(clk),
	.Q(currMEM[31]));
   DFF_X1 currMEM_reg_30_ (.D(n98),
	.CK(clk),
	.Q(currMEM[30]));
   DFF_X1 currMEM_reg_29_ (.D(n99),
	.CK(clk),
	.Q(currMEM[29]));
   DFF_X1 currMEM_reg_28_ (.D(n100),
	.CK(clk),
	.Q(currMEM[28]));
   DFF_X1 currMEM_reg_27_ (.D(n101),
	.CK(clk),
	.Q(currMEM[27]));
   DFF_X1 currMEM_reg_26_ (.D(n102),
	.CK(clk),
	.Q(currMEM[26]));
   DFF_X1 currMEM_reg_25_ (.D(n206),
	.CK(clk),
	.Q(currMEM[25]));
   DFF_X1 currMEM_reg_24_ (.D(n207),
	.CK(clk),
	.Q(currMEM[24]));
   DFF_X1 currMEM_reg_23_ (.D(n208),
	.CK(clk),
	.Q(currMEM[23]));
   DFF_X1 currMEM_reg_22_ (.D(n209),
	.CK(clk),
	.Q(currMEM[22]));
   DFF_X1 currMEM_reg_21_ (.D(n210),
	.CK(clk),
	.Q(currMEM[21]));
   DFF_X1 currMEM_reg_20_ (.D(n211),
	.CK(clk),
	.Q(currMEM[20]));
   DFF_X1 currMEM_reg_19_ (.D(n212),
	.CK(clk),
	.Q(currMEM[19]));
   DFF_X1 currMEM_reg_18_ (.D(n213),
	.CK(clk),
	.Q(currMEM[18]));
   DFF_X1 currMEM_reg_17_ (.D(n214),
	.CK(clk),
	.Q(currMEM[17]));
   DFF_X1 currMEM_reg_16_ (.D(n215),
	.CK(clk),
	.Q(currMEM[16]));
   DFF_X1 currMEM_reg_15_ (.D(n216),
	.CK(clk),
	.Q(currMEM[15]));
   DFF_X1 currMEM_reg_14_ (.D(n217),
	.CK(clk),
	.Q(currMEM[14]));
   DFF_X1 currMEM_reg_13_ (.D(n218),
	.CK(clk),
	.Q(currMEM[13]));
   DFF_X1 currMEM_reg_12_ (.D(n219),
	.CK(clk),
	.Q(currMEM[12]));
   DFF_X1 currMEM_reg_11_ (.D(n220),
	.CK(clk),
	.Q(currMEM[11]));
   DFF_X1 currMEM_reg_10_ (.D(n221),
	.CK(clk),
	.Q(currMEM[10]));
   DFF_X1 currMEM_reg_9_ (.D(n222),
	.CK(clk),
	.Q(currMEM[9]));
   DFF_X1 currMEM_reg_8_ (.D(n223),
	.CK(clk),
	.Q(currMEM[8]));
   DFF_X1 currMEM_reg_7_ (.D(n224),
	.CK(clk),
	.Q(currMEM[7]));
   DFF_X1 currMEM_reg_6_ (.D(n225),
	.CK(clk),
	.Q(currMEM[6]));
   DFF_X1 currMEM_reg_5_ (.D(n226),
	.CK(clk),
	.Q(currMEM[5]));
   DFF_X1 currMEM_reg_4_ (.D(n227),
	.CK(clk),
	.Q(currMEM[4]));
   DFF_X1 currMEM_reg_3_ (.D(n228),
	.CK(clk),
	.Q(currMEM[3]));
   DFF_X1 currMEM_reg_2_ (.D(n229),
	.CK(clk),
	.Q(currMEM[2]));
   DFF_X1 currMEM_reg_1_ (.D(n230),
	.CK(clk),
	.Q(currMEM[1]));
   DFF_X1 currMEM_reg_0_ (.D(n231),
	.CK(clk),
	.Q(currMEM[0]));
   DFF_X1 currRD_reg_0_ (.D(n32),
	.CK(clk),
	.Q(RD_OUT[0]),
	.QN(n3));
   DFF_X1 currRD_reg_1_ (.D(n31),
	.CK(clk),
	.Q(RD_OUT[1]));
   DFF_X1 currRD_reg_2_ (.D(n30),
	.CK(clk),
	.Q(RD_OUT[2]),
	.QN(n1));
   DFF_X2 currRD_reg_4_ (.D(n28),
	.CK(clk),
	.Q(RD_OUT[4]));
   DFF_X1 currRD_reg_3_ (.D(n29),
	.CK(clk),
	.Q(RD_OUT[3]));
   INV_X1 U3 (.A(n1),
	.ZN(n2));
   INV_X1 U4 (.A(n3),
	.ZN(n4));
   INV_X2 U5 (.A(MUX_SEL),
	.ZN(n27));
   INV_X1 U27 (.A(n202),
	.ZN(WB_OUT[12]));
   AOI22_X1 U28 (.A1(currMEM[12]),
	.A2(MUX_SEL),
	.B1(n27),
	.B2(currALU[12]),
	.ZN(n202));
   INV_X1 U29 (.A(n183),
	.ZN(WB_OUT[2]));
   AOI22_X1 U30 (.A1(currMEM[2]),
	.A2(FE_OFN41_MUX_SEL_WB_c),
	.B1(n27),
	.B2(currALU[2]),
	.ZN(n183));
   INV_X1 U31 (.A(n175),
	.ZN(WB_OUT[8]));
   AOI22_X1 U32 (.A1(currMEM[8]),
	.A2(MUX_SEL),
	.B1(n27),
	.B2(currALU[8]),
	.ZN(n175));
   INV_X1 U33 (.A(n180),
	.ZN(WB_OUT[3]));
   AOI22_X1 U34 (.A1(currMEM[3]),
	.A2(FE_OFN41_MUX_SEL_WB_c),
	.B1(n27),
	.B2(currALU[3]),
	.ZN(n180));
   INV_X1 U35 (.A(n179),
	.ZN(WB_OUT[4]));
   AOI22_X1 U36 (.A1(currMEM[4]),
	.A2(MUX_SEL),
	.B1(n27),
	.B2(currALU[4]),
	.ZN(n179));
   INV_X1 U37 (.A(n174),
	.ZN(WB_OUT[9]));
   AOI22_X1 U38 (.A1(currMEM[9]),
	.A2(MUX_SEL),
	.B1(n27),
	.B2(currALU[9]),
	.ZN(n174));
   INV_X1 U39 (.A(n178),
	.ZN(WB_OUT[5]));
   AOI22_X1 U40 (.A1(currMEM[5]),
	.A2(MUX_SEL),
	.B1(n27),
	.B2(currALU[5]),
	.ZN(n178));
   INV_X1 U41 (.A(n177),
	.ZN(WB_OUT[6]));
   AOI22_X1 U42 (.A1(currMEM[6]),
	.A2(FE_OFN41_MUX_SEL_WB_c),
	.B1(n27),
	.B2(currALU[6]),
	.ZN(n177));
   INV_X1 U43 (.A(n176),
	.ZN(WB_OUT[7]));
   AOI22_X1 U44 (.A1(currMEM[7]),
	.A2(MUX_SEL),
	.B1(n27),
	.B2(currALU[7]),
	.ZN(n176));
   INV_X1 U45 (.A(n205),
	.ZN(WB_OUT[0]));
   AOI22_X1 U46 (.A1(currMEM[0]),
	.A2(MUX_SEL),
	.B1(n27),
	.B2(currALU[0]),
	.ZN(n205));
   INV_X1 U47 (.A(n194),
	.ZN(WB_OUT[1]));
   AOI22_X1 U48 (.A1(currMEM[1]),
	.A2(FE_OFN41_MUX_SEL_WB_c),
	.B1(n27),
	.B2(currALU[1]),
	.ZN(n194));
   INV_X1 U49 (.A(n204),
	.ZN(WB_OUT[10]));
   AOI22_X1 U50 (.A1(currMEM[10]),
	.A2(MUX_SEL),
	.B1(n27),
	.B2(currALU[10]),
	.ZN(n204));
   INV_X1 U51 (.A(n203),
	.ZN(WB_OUT[11]));
   AOI22_X1 U52 (.A1(currMEM[11]),
	.A2(MUX_SEL),
	.B1(n27),
	.B2(currALU[11]),
	.ZN(n203));
   INV_X1 U53 (.A(n201),
	.ZN(WB_OUT[13]));
   AOI22_X1 U54 (.A1(currMEM[13]),
	.A2(FE_OFN41_MUX_SEL_WB_c),
	.B1(n27),
	.B2(currALU[13]),
	.ZN(n201));
   INV_X1 U55 (.A(n200),
	.ZN(WB_OUT[14]));
   AOI22_X1 U56 (.A1(currMEM[14]),
	.A2(MUX_SEL),
	.B1(n27),
	.B2(currALU[14]),
	.ZN(n200));
   INV_X1 U57 (.A(n199),
	.ZN(WB_OUT[15]));
   AOI22_X1 U58 (.A1(currMEM[15]),
	.A2(MUX_SEL),
	.B1(n27),
	.B2(currALU[15]),
	.ZN(n199));
   INV_X1 U59 (.A(n198),
	.ZN(WB_OUT[16]));
   AOI22_X1 U60 (.A1(currMEM[16]),
	.A2(MUX_SEL),
	.B1(n27),
	.B2(currALU[16]),
	.ZN(n198));
   INV_X1 U61 (.A(n197),
	.ZN(WB_OUT[17]));
   AOI22_X1 U62 (.A1(currMEM[17]),
	.A2(FE_OFN41_MUX_SEL_WB_c),
	.B1(n27),
	.B2(currALU[17]),
	.ZN(n197));
   INV_X1 U63 (.A(n196),
	.ZN(WB_OUT[18]));
   AOI22_X1 U64 (.A1(currMEM[18]),
	.A2(FE_OFN41_MUX_SEL_WB_c),
	.B1(n27),
	.B2(currALU[18]),
	.ZN(n196));
   INV_X1 U65 (.A(n181),
	.ZN(WB_OUT[31]));
   AOI22_X1 U66 (.A1(currMEM[31]),
	.A2(FE_OFN41_MUX_SEL_WB_c),
	.B1(n27),
	.B2(currALU[31]),
	.ZN(n181));
   INV_X1 U67 (.A(n182),
	.ZN(WB_OUT[30]));
   AOI22_X1 U68 (.A1(currMEM[30]),
	.A2(FE_OFN41_MUX_SEL_WB_c),
	.B1(n27),
	.B2(currALU[30]),
	.ZN(n182));
   INV_X1 U69 (.A(n184),
	.ZN(WB_OUT[29]));
   AOI22_X1 U70 (.A1(currMEM[29]),
	.A2(FE_OFN41_MUX_SEL_WB_c),
	.B1(n27),
	.B2(currALU[29]),
	.ZN(n184));
   INV_X1 U71 (.A(n193),
	.ZN(WB_OUT[20]));
   AOI22_X1 U72 (.A1(currMEM[20]),
	.A2(FE_OFN41_MUX_SEL_WB_c),
	.B1(n27),
	.B2(currALU[20]),
	.ZN(n193));
   INV_X1 U73 (.A(n192),
	.ZN(WB_OUT[21]));
   AOI22_X1 U74 (.A1(currMEM[21]),
	.A2(FE_OFN41_MUX_SEL_WB_c),
	.B1(n27),
	.B2(currALU[21]),
	.ZN(n192));
   INV_X1 U75 (.A(n191),
	.ZN(WB_OUT[22]));
   AOI22_X1 U76 (.A1(currMEM[22]),
	.A2(FE_OFN41_MUX_SEL_WB_c),
	.B1(n27),
	.B2(currALU[22]),
	.ZN(n191));
   INV_X1 U77 (.A(n190),
	.ZN(WB_OUT[23]));
   AOI22_X1 U78 (.A1(currMEM[23]),
	.A2(FE_OFN41_MUX_SEL_WB_c),
	.B1(n27),
	.B2(currALU[23]),
	.ZN(n190));
   INV_X1 U79 (.A(n189),
	.ZN(WB_OUT[24]));
   AOI22_X1 U80 (.A1(currMEM[24]),
	.A2(FE_OFN41_MUX_SEL_WB_c),
	.B1(n27),
	.B2(currALU[24]),
	.ZN(n189));
   INV_X1 U81 (.A(n188),
	.ZN(WB_OUT[25]));
   AOI22_X1 U82 (.A1(currMEM[25]),
	.A2(FE_OFN41_MUX_SEL_WB_c),
	.B1(n27),
	.B2(currALU[25]),
	.ZN(n188));
   INV_X1 U83 (.A(n187),
	.ZN(WB_OUT[26]));
   AOI22_X1 U84 (.A1(currMEM[26]),
	.A2(FE_OFN41_MUX_SEL_WB_c),
	.B1(n27),
	.B2(currALU[26]),
	.ZN(n187));
   INV_X1 U85 (.A(n186),
	.ZN(WB_OUT[27]));
   AOI22_X1 U86 (.A1(currMEM[27]),
	.A2(FE_OFN41_MUX_SEL_WB_c),
	.B1(n27),
	.B2(currALU[27]),
	.ZN(n186));
   INV_X1 U87 (.A(n185),
	.ZN(WB_OUT[28]));
   AOI22_X1 U88 (.A1(currMEM[28]),
	.A2(FE_OFN41_MUX_SEL_WB_c),
	.B1(n27),
	.B2(currALU[28]),
	.ZN(n185));
   INV_X1 U89 (.A(n195),
	.ZN(WB_OUT[19]));
   AOI22_X1 U90 (.A1(currMEM[19]),
	.A2(FE_OFN41_MUX_SEL_WB_c),
	.B1(n27),
	.B2(currALU[19]),
	.ZN(n195));
   NOR2_X1 U91 (.A1(en),
	.A2(rst),
	.ZN(n104));
   NOR2_X1 U92 (.A1(FE_OFN15_n104),
	.A2(rst),
	.ZN(n105));
   INV_X1 U93 (.A(n171),
	.ZN(n30));
   INV_X1 U94 (.A(n170),
	.ZN(n31));
   INV_X1 U95 (.A(n173),
	.ZN(n28));
   AOI22_X1 U96 (.A1(RD_IN[4]),
	.A2(n105),
	.B1(RD_OUT[4]),
	.B2(n104),
	.ZN(n173));
   INV_X1 U97 (.A(n172),
	.ZN(n29));
   AOI22_X1 U98 (.A1(RD_IN[3]),
	.A2(n105),
	.B1(RD_OUT[3]),
	.B2(n104),
	.ZN(n172));
   INV_X1 U99 (.A(n169),
	.ZN(n32));
   INV_X1 U100 (.A(n162),
	.ZN(n46));
   AOI22_X1 U101 (.A1(FE_OFN15_n104),
	.A2(currALU[25]),
	.B1(FE_OFN57_n105),
	.B2(ALU_OUT[25]),
	.ZN(n162));
   INV_X1 U102 (.A(n163),
	.ZN(n44));
   AOI22_X1 U103 (.A1(FE_OFN16_n104),
	.A2(currALU[26]),
	.B1(FE_OFN57_n105),
	.B2(ALU_OUT[26]),
	.ZN(n163));
   INV_X1 U104 (.A(n164),
	.ZN(n42));
   AOI22_X1 U105 (.A1(FE_OFN15_n104),
	.A2(currALU[27]),
	.B1(FE_OFN57_n105),
	.B2(ALU_OUT[27]),
	.ZN(n164));
   INV_X1 U106 (.A(n165),
	.ZN(n40));
   AOI22_X1 U107 (.A1(FE_OFN16_n104),
	.A2(currALU[28]),
	.B1(FE_OFN57_n105),
	.B2(ALU_OUT[28]),
	.ZN(n165));
   INV_X1 U108 (.A(n166),
	.ZN(n38));
   AOI22_X1 U109 (.A1(FE_OFN16_n104),
	.A2(currALU[29]),
	.B1(FE_OFN57_n105),
	.B2(ALU_OUT[29]),
	.ZN(n166));
   INV_X1 U110 (.A(n167),
	.ZN(n36));
   AOI22_X1 U111 (.A1(FE_OFN16_n104),
	.A2(currALU[30]),
	.B1(FE_OFN57_n105),
	.B2(ALU_OUT[30]),
	.ZN(n167));
   INV_X1 U112 (.A(n139),
	.ZN(n92));
   AOI22_X1 U113 (.A1(FE_OFN15_n104),
	.A2(currALU[2]),
	.B1(FE_OFN57_n105),
	.B2(ALU_OUT[2]),
	.ZN(n139));
   INV_X1 U114 (.A(n103),
	.ZN(n231));
   AOI22_X1 U115 (.A1(FE_OFN15_n104),
	.A2(currMEM[0]),
	.B1(FE_OFN57_n105),
	.B2(DRAM_OUT[0]),
	.ZN(n103));
   INV_X1 U116 (.A(n137),
	.ZN(n96));
   AOI22_X1 U117 (.A1(FE_OFN15_n104),
	.A2(currALU[0]),
	.B1(FE_OFN57_n105),
	.B2(ALU_OUT[0]),
	.ZN(n137));
   INV_X1 U118 (.A(n138),
	.ZN(n94));
   AOI22_X1 U119 (.A1(FE_OFN15_n104),
	.A2(currALU[1]),
	.B1(FE_OFN57_n105),
	.B2(ALU_OUT[1]),
	.ZN(n138));
   INV_X1 U120 (.A(n140),
	.ZN(n90));
   AOI22_X1 U121 (.A1(FE_OFN15_n104),
	.A2(currALU[3]),
	.B1(FE_OFN57_n105),
	.B2(ALU_OUT[3]),
	.ZN(n140));
   INV_X1 U122 (.A(n141),
	.ZN(n88));
   AOI22_X1 U123 (.A1(FE_OFN15_n104),
	.A2(currALU[4]),
	.B1(FE_OFN57_n105),
	.B2(ALU_OUT[4]),
	.ZN(n141));
   INV_X1 U124 (.A(n142),
	.ZN(n86));
   AOI22_X1 U125 (.A1(FE_OFN15_n104),
	.A2(currALU[5]),
	.B1(FE_OFN57_n105),
	.B2(ALU_OUT[5]),
	.ZN(n142));
   INV_X1 U126 (.A(n143),
	.ZN(n84));
   AOI22_X1 U127 (.A1(FE_OFN15_n104),
	.A2(currALU[6]),
	.B1(FE_OFN57_n105),
	.B2(ALU_OUT[6]),
	.ZN(n143));
   INV_X1 U128 (.A(n144),
	.ZN(n82));
   AOI22_X1 U129 (.A1(FE_OFN15_n104),
	.A2(currALU[7]),
	.B1(FE_OFN57_n105),
	.B2(ALU_OUT[7]),
	.ZN(n144));
   INV_X1 U130 (.A(n145),
	.ZN(n80));
   AOI22_X1 U131 (.A1(FE_OFN15_n104),
	.A2(currALU[8]),
	.B1(FE_OFN57_n105),
	.B2(ALU_OUT[8]),
	.ZN(n145));
   INV_X1 U132 (.A(n146),
	.ZN(n78));
   AOI22_X1 U133 (.A1(FE_OFN15_n104),
	.A2(currALU[9]),
	.B1(FE_OFN57_n105),
	.B2(ALU_OUT[9]),
	.ZN(n146));
   INV_X1 U134 (.A(n147),
	.ZN(n76));
   AOI22_X1 U135 (.A1(FE_OFN15_n104),
	.A2(currALU[10]),
	.B1(FE_OFN57_n105),
	.B2(ALU_OUT[10]),
	.ZN(n147));
   INV_X1 U136 (.A(n148),
	.ZN(n74));
   AOI22_X1 U137 (.A1(FE_OFN15_n104),
	.A2(currALU[11]),
	.B1(FE_OFN57_n105),
	.B2(ALU_OUT[11]),
	.ZN(n148));
   INV_X1 U138 (.A(n149),
	.ZN(n72));
   AOI22_X1 U139 (.A1(FE_OFN15_n104),
	.A2(currALU[12]),
	.B1(FE_OFN57_n105),
	.B2(ALU_OUT[12]),
	.ZN(n149));
   INV_X1 U140 (.A(n150),
	.ZN(n70));
   AOI22_X1 U141 (.A1(FE_OFN15_n104),
	.A2(currALU[13]),
	.B1(FE_OFN57_n105),
	.B2(ALU_OUT[13]),
	.ZN(n150));
   INV_X1 U142 (.A(n151),
	.ZN(n68));
   AOI22_X1 U143 (.A1(FE_OFN15_n104),
	.A2(currALU[14]),
	.B1(FE_OFN57_n105),
	.B2(ALU_OUT[14]),
	.ZN(n151));
   INV_X1 U144 (.A(n152),
	.ZN(n66));
   AOI22_X1 U145 (.A1(FE_OFN15_n104),
	.A2(currALU[15]),
	.B1(FE_OFN57_n105),
	.B2(ALU_OUT[15]),
	.ZN(n152));
   INV_X1 U146 (.A(n153),
	.ZN(n64));
   AOI22_X1 U147 (.A1(FE_OFN15_n104),
	.A2(currALU[16]),
	.B1(FE_OFN57_n105),
	.B2(ALU_OUT[16]),
	.ZN(n153));
   INV_X1 U148 (.A(n154),
	.ZN(n62));
   AOI22_X1 U149 (.A1(FE_OFN15_n104),
	.A2(currALU[17]),
	.B1(FE_OFN57_n105),
	.B2(ALU_OUT[17]),
	.ZN(n154));
   INV_X1 U150 (.A(n155),
	.ZN(n60));
   AOI22_X1 U151 (.A1(FE_OFN16_n104),
	.A2(currALU[18]),
	.B1(FE_OFN57_n105),
	.B2(ALU_OUT[18]),
	.ZN(n155));
   INV_X1 U152 (.A(n156),
	.ZN(n58));
   AOI22_X1 U153 (.A1(FE_OFN15_n104),
	.A2(currALU[19]),
	.B1(FE_OFN57_n105),
	.B2(ALU_OUT[19]),
	.ZN(n156));
   INV_X1 U154 (.A(n157),
	.ZN(n56));
   AOI22_X1 U155 (.A1(FE_OFN16_n104),
	.A2(currALU[20]),
	.B1(FE_OFN57_n105),
	.B2(ALU_OUT[20]),
	.ZN(n157));
   INV_X1 U156 (.A(n158),
	.ZN(n54));
   AOI22_X1 U157 (.A1(FE_OFN16_n104),
	.A2(currALU[21]),
	.B1(FE_OFN57_n105),
	.B2(ALU_OUT[21]),
	.ZN(n158));
   INV_X1 U158 (.A(n159),
	.ZN(n52));
   AOI22_X1 U159 (.A1(FE_OFN16_n104),
	.A2(currALU[22]),
	.B1(FE_OFN57_n105),
	.B2(ALU_OUT[22]),
	.ZN(n159));
   INV_X1 U160 (.A(n160),
	.ZN(n50));
   AOI22_X1 U161 (.A1(FE_OFN16_n104),
	.A2(currALU[23]),
	.B1(FE_OFN57_n105),
	.B2(ALU_OUT[23]),
	.ZN(n160));
   INV_X1 U162 (.A(n161),
	.ZN(n48));
   AOI22_X1 U163 (.A1(FE_OFN16_n104),
	.A2(currALU[24]),
	.B1(FE_OFN57_n105),
	.B2(ALU_OUT[24]),
	.ZN(n161));
   INV_X1 U164 (.A(n106),
	.ZN(n230));
   AOI22_X1 U165 (.A1(FE_OFN15_n104),
	.A2(currMEM[1]),
	.B1(FE_OFN57_n105),
	.B2(DRAM_OUT[1]),
	.ZN(n106));
   INV_X1 U166 (.A(n107),
	.ZN(n229));
   AOI22_X1 U167 (.A1(FE_OFN15_n104),
	.A2(currMEM[2]),
	.B1(FE_OFN57_n105),
	.B2(DRAM_OUT[2]),
	.ZN(n107));
   INV_X1 U168 (.A(n108),
	.ZN(n228));
   AOI22_X1 U169 (.A1(FE_OFN15_n104),
	.A2(currMEM[3]),
	.B1(FE_OFN57_n105),
	.B2(DRAM_OUT[3]),
	.ZN(n108));
   INV_X1 U170 (.A(n109),
	.ZN(n227));
   AOI22_X1 U171 (.A1(FE_OFN15_n104),
	.A2(currMEM[4]),
	.B1(n105),
	.B2(DRAM_OUT[4]),
	.ZN(n109));
   INV_X1 U172 (.A(n110),
	.ZN(n226));
   AOI22_X1 U173 (.A1(FE_OFN15_n104),
	.A2(currMEM[5]),
	.B1(FE_OFN57_n105),
	.B2(DRAM_OUT[5]),
	.ZN(n110));
   INV_X1 U174 (.A(n111),
	.ZN(n225));
   AOI22_X1 U175 (.A1(FE_OFN15_n104),
	.A2(currMEM[6]),
	.B1(FE_OFN57_n105),
	.B2(DRAM_OUT[6]),
	.ZN(n111));
   INV_X1 U176 (.A(n112),
	.ZN(n224));
   AOI22_X1 U177 (.A1(FE_OFN15_n104),
	.A2(currMEM[7]),
	.B1(FE_OFN57_n105),
	.B2(DRAM_OUT[7]),
	.ZN(n112));
   INV_X1 U178 (.A(n113),
	.ZN(n223));
   AOI22_X1 U179 (.A1(FE_OFN15_n104),
	.A2(currMEM[8]),
	.B1(FE_OFN57_n105),
	.B2(DRAM_OUT[8]),
	.ZN(n113));
   INV_X1 U180 (.A(n114),
	.ZN(n222));
   AOI22_X1 U181 (.A1(FE_OFN15_n104),
	.A2(currMEM[9]),
	.B1(FE_OFN57_n105),
	.B2(DRAM_OUT[9]),
	.ZN(n114));
   INV_X1 U182 (.A(n115),
	.ZN(n221));
   AOI22_X1 U183 (.A1(FE_OFN15_n104),
	.A2(currMEM[10]),
	.B1(FE_OFN57_n105),
	.B2(DRAM_OUT[10]),
	.ZN(n115));
   INV_X1 U184 (.A(n116),
	.ZN(n220));
   AOI22_X1 U185 (.A1(FE_OFN15_n104),
	.A2(currMEM[11]),
	.B1(n105),
	.B2(DRAM_OUT[11]),
	.ZN(n116));
   INV_X1 U186 (.A(n117),
	.ZN(n219));
   AOI22_X1 U187 (.A1(FE_OFN15_n104),
	.A2(currMEM[12]),
	.B1(FE_OFN57_n105),
	.B2(DRAM_OUT[12]),
	.ZN(n117));
   INV_X1 U188 (.A(n118),
	.ZN(n218));
   AOI22_X1 U189 (.A1(FE_OFN15_n104),
	.A2(currMEM[13]),
	.B1(FE_OFN57_n105),
	.B2(DRAM_OUT[13]),
	.ZN(n118));
   INV_X1 U190 (.A(n119),
	.ZN(n217));
   AOI22_X1 U191 (.A1(FE_OFN15_n104),
	.A2(currMEM[14]),
	.B1(FE_OFN57_n105),
	.B2(DRAM_OUT[14]),
	.ZN(n119));
   INV_X1 U192 (.A(n120),
	.ZN(n216));
   AOI22_X1 U193 (.A1(FE_OFN15_n104),
	.A2(currMEM[15]),
	.B1(FE_OFN57_n105),
	.B2(DRAM_OUT[15]),
	.ZN(n120));
   INV_X1 U194 (.A(n121),
	.ZN(n215));
   AOI22_X1 U195 (.A1(FE_OFN15_n104),
	.A2(currMEM[16]),
	.B1(FE_OFN57_n105),
	.B2(DRAM_OUT[16]),
	.ZN(n121));
   INV_X1 U196 (.A(n122),
	.ZN(n214));
   AOI22_X1 U197 (.A1(FE_OFN15_n104),
	.A2(currMEM[17]),
	.B1(FE_OFN57_n105),
	.B2(DRAM_OUT[17]),
	.ZN(n122));
   INV_X1 U198 (.A(n123),
	.ZN(n213));
   AOI22_X1 U199 (.A1(FE_OFN16_n104),
	.A2(currMEM[18]),
	.B1(FE_OFN57_n105),
	.B2(DRAM_OUT[18]),
	.ZN(n123));
   INV_X1 U200 (.A(n124),
	.ZN(n212));
   AOI22_X1 U201 (.A1(FE_OFN15_n104),
	.A2(currMEM[19]),
	.B1(FE_OFN57_n105),
	.B2(DRAM_OUT[19]),
	.ZN(n124));
   INV_X1 U202 (.A(n125),
	.ZN(n211));
   AOI22_X1 U203 (.A1(FE_OFN16_n104),
	.A2(currMEM[20]),
	.B1(FE_OFN57_n105),
	.B2(DRAM_OUT[20]),
	.ZN(n125));
   INV_X1 U204 (.A(n126),
	.ZN(n210));
   AOI22_X1 U205 (.A1(FE_OFN16_n104),
	.A2(currMEM[21]),
	.B1(FE_OFN57_n105),
	.B2(DRAM_OUT[21]),
	.ZN(n126));
   INV_X1 U206 (.A(n127),
	.ZN(n209));
   AOI22_X1 U207 (.A1(FE_OFN16_n104),
	.A2(currMEM[22]),
	.B1(FE_OFN57_n105),
	.B2(DRAM_OUT[22]),
	.ZN(n127));
   INV_X1 U208 (.A(n128),
	.ZN(n208));
   AOI22_X1 U209 (.A1(FE_OFN16_n104),
	.A2(currMEM[23]),
	.B1(FE_OFN57_n105),
	.B2(DRAM_OUT[23]),
	.ZN(n128));
   INV_X1 U210 (.A(n129),
	.ZN(n207));
   AOI22_X1 U211 (.A1(FE_OFN16_n104),
	.A2(currMEM[24]),
	.B1(FE_OFN57_n105),
	.B2(DRAM_OUT[24]),
	.ZN(n129));
   INV_X1 U212 (.A(n130),
	.ZN(n206));
   AOI22_X1 U213 (.A1(FE_OFN15_n104),
	.A2(currMEM[25]),
	.B1(FE_OFN57_n105),
	.B2(DRAM_OUT[25]),
	.ZN(n130));
   INV_X1 U214 (.A(n131),
	.ZN(n102));
   AOI22_X1 U215 (.A1(FE_OFN16_n104),
	.A2(currMEM[26]),
	.B1(FE_OFN57_n105),
	.B2(DRAM_OUT[26]),
	.ZN(n131));
   INV_X1 U216 (.A(n132),
	.ZN(n101));
   AOI22_X1 U217 (.A1(FE_OFN15_n104),
	.A2(currMEM[27]),
	.B1(FE_OFN57_n105),
	.B2(DRAM_OUT[27]),
	.ZN(n132));
   INV_X1 U218 (.A(n133),
	.ZN(n100));
   AOI22_X1 U219 (.A1(FE_OFN16_n104),
	.A2(currMEM[28]),
	.B1(FE_OFN57_n105),
	.B2(DRAM_OUT[28]),
	.ZN(n133));
   INV_X1 U220 (.A(n134),
	.ZN(n99));
   AOI22_X1 U221 (.A1(FE_OFN16_n104),
	.A2(currMEM[29]),
	.B1(FE_OFN57_n105),
	.B2(DRAM_OUT[29]),
	.ZN(n134));
   INV_X1 U222 (.A(n135),
	.ZN(n98));
   AOI22_X1 U223 (.A1(FE_OFN16_n104),
	.A2(currMEM[30]),
	.B1(FE_OFN57_n105),
	.B2(DRAM_OUT[30]),
	.ZN(n135));
   INV_X1 U224 (.A(n136),
	.ZN(n97));
   AOI22_X1 U225 (.A1(FE_OFN16_n104),
	.A2(currMEM[31]),
	.B1(FE_OFN57_n105),
	.B2(DRAM_OUT[31]),
	.ZN(n136));
   INV_X1 U226 (.A(n168),
	.ZN(n34));
   AOI22_X1 U227 (.A1(FE_OFN16_n104),
	.A2(currALU[31]),
	.B1(FE_OFN57_n105),
	.B2(ALU_OUT[31]),
	.ZN(n168));
   AOI22_X1 U228 (.A1(RD_IN[2]),
	.A2(n105),
	.B1(n2),
	.B2(n104),
	.ZN(n171));
   AOI22_X1 U229 (.A1(RD_IN[1]),
	.A2(n105),
	.B1(RD_OUT[1]),
	.B2(n104),
	.ZN(n170));
   AOI22_X1 U230 (.A1(RD_IN[0]),
	.A2(n105),
	.B1(n4),
	.B2(n104),
	.ZN(n169));
endmodule

module DP (
	clk, 
	rst, 
	FETCH_EN, 
	DECODE_EN, 
	EXE_EN, 
	MEM_EN, 
	WB_EN, 
	IRAM_OUT, 
	DRAM_OUT, 
	DRAM_WR_IN, 
	DRAM_RD_IN, 
	RF_RD1, 
	RF_RD2, 
	RF_WR, 
	JUMP, 
	MUX_SEL_WB, 
	RF_OUT1_SEL, 
	RF_OUT2_SEL, 
	ALU_OPA_SEL, 
	ALU_OPB_SEL, 
	MUX_SEL_IMM, 
	ALU_OP, 
	IRAM_ADDR, 
	DRAM_IN, 
	DRAM_ADDR, 
	DRAM_WR, 
	DRAM_RD, 
	OPCODE, 
	FUNC3, 
	EQU, 
	RS1_IF_ID, 
	RS2_IF_ID, 
	RS1_ID_EXE, 
	RS2_ID_EXE, 
	RD_EXE_MEM, 
	RD_MEM_WB, 
	RD_ID_EXE);
   input clk;
   input rst;
   input FETCH_EN;
   input DECODE_EN;
   input EXE_EN;
   input MEM_EN;
   input WB_EN;
   input [31:0] IRAM_OUT;
   input [31:0] DRAM_OUT;
   input DRAM_WR_IN;
   input DRAM_RD_IN;
   input RF_RD1;
   input RF_RD2;
   input RF_WR;
   input JUMP;
   input MUX_SEL_WB;
   input [1:0] RF_OUT1_SEL;
   input [1:0] RF_OUT2_SEL;
   input [2:0] ALU_OPA_SEL;
   input [2:0] ALU_OPB_SEL;
   input [2:0] MUX_SEL_IMM;
   input [2:0] ALU_OP;
   output [31:0] IRAM_ADDR;
   output [31:0] DRAM_IN;
   output [31:0] DRAM_ADDR;
   output DRAM_WR;
   output DRAM_RD;
   output [6:0] OPCODE;
   output [2:0] FUNC3;
   output EQU;
   output [4:0] RS1_IF_ID;
   output [4:0] RS2_IF_ID;
   output [4:0] RS1_ID_EXE;
   output [4:0] RS2_ID_EXE;
   output [4:0] RD_EXE_MEM;
   output [4:0] RD_MEM_WB;
   output [4:0] RD_ID_EXE;

   // Internal wires
   wire [31:0] pc_jump_addr_m;
   wire [31:0] ir_m;
   wire [31:0] wb_out_m;
   wire [31:0] rf_out1_m;
   wire [31:0] rf_out2_m;
   wire [31:0] pc_ext_m;
   wire [31:0] imm_m;
   wire [4:0] rd_m1;
   wire [31:0] alu_out_m1;
   wire [31:0] mem_data_m;
   wire [31:0] dram_out_m;

   fetch_unit FETCH_U (.clk(clk),
	.rst(rst),
	.en(FETCH_EN),
	.PC_MUX_SEL(JUMP),
	.IRAM_DOUT_IN(IRAM_OUT),
	.PC_JUMP_ADDR(pc_jump_addr_m),
	.PC(IRAM_ADDR),
	.IR_IN(ir_m));
   decode_unit DECODE_U (.clk(clk),
	.rst(rst),
	.en(DECODE_EN),
	.RF_RD1(RF_RD1),
	.RF_RD2(RF_RD2),
	.RF_WR(RF_WR),
	.IF_FLUSH(JUMP),
	.PC_IN(IRAM_ADDR),
	.IR_IN(ir_m),
	.EXE_MEM_IN(DRAM_ADDR),
	.ADD_WR(RD_MEM_WB),
	.DATAIN(wb_out_m),
	.MUX_IMM_SEL(MUX_SEL_IMM),
	.RF_OUT1_SEL(RF_OUT1_SEL),
	.RF_OUT2_SEL(RF_OUT2_SEL),
	.OPCODE(OPCODE),
	.FUNC3(FUNC3),
	.EQU_FLAG(EQU),
	.RF_OUT1(rf_out1_m),
	.RF_OUT2(rf_out2_m),
	.PC_OUT(pc_ext_m),
	.IMM(imm_m),
	.JMP_ADDR(pc_jump_addr_m),
	.RD(rd_m1),
	.RS1(RS1_IF_ID),
	.RS2(RS2_IF_ID));
   exe_unit EXE_U (.clk(clk),
	.rst(rst),
	.en(EXE_EN),
	.RF_OUT1(rf_out1_m),
	.RF_OUT2(rf_out2_m),
	.PC(pc_ext_m),
	.IMM(imm_m),
	.EXE_MEM_IN(DRAM_ADDR),
	.MEM_WB_IN(wb_out_m),
	.RD_IN(rd_m1),
	.RS1_IN(RS1_IF_ID),
	.RS2_IN(RS2_IF_ID),
	.ALU_OP(ALU_OP),
	.ALU_OPA_SEL(ALU_OPA_SEL),
	.ALU_OPB_SEL(ALU_OPB_SEL),
	.ALU_OUT(alu_out_m1),
	.MEM_DATA(mem_data_m),
	.RD_OUT(RD_ID_EXE),
	.RS1_OUT(RS1_ID_EXE),
	.RS2_OUT(RS2_ID_EXE));
   mem_unit MEM_U (.clk(clk),
	.rst(rst),
	.en(MEM_EN),
	.ALU_OUT_IN(alu_out_m1),
	.MEM_DATA(mem_data_m),
	.DRAM_OUT_IN(DRAM_OUT),
	.DRAM_WR_IN(DRAM_WR_IN),
	.DRAM_RD_IN(DRAM_RD_IN),
	.RD_IN(RD_ID_EXE),
	.RD_OUT(RD_EXE_MEM),
	.DRAM_WR(DRAM_WR),
	.DRAM_RD(DRAM_RD),
	.ALU_OUT(DRAM_ADDR),
	.DRAM_OUT(dram_out_m),
	.DRAM_IN(DRAM_IN));
   wb_unit WB_U (.clk(clk),
	.rst(rst),
	.en(WB_EN),
	.RD_IN(RD_EXE_MEM),
	.ALU_OUT(DRAM_ADDR),
	.DRAM_OUT(dram_out_m),
	.MUX_SEL(MUX_SEL_WB),
	.RD_OUT(RD_MEM_WB),
	.WB_OUT(wb_out_m));
endmodule

module FWD_EXE (
	RS1_ID_EX, 
	RS2_ID_EX, 
	RD_EX_MEM, 
	RD_MEM_WB, 
	MUX_OPA_SEL_STD, 
	MUX_OPB_SEL_STD, 
	EXE_MEM_WR, 
	MEM_WB_WR, 
	MUX_OPA_SEL, 
	MUX_OPB_SEL);
   input [4:0] RS1_ID_EX;
   input [4:0] RS2_ID_EX;
   input [4:0] RD_EX_MEM;
   input [4:0] RD_MEM_WB;
   input [2:0] MUX_OPA_SEL_STD;
   input [2:0] MUX_OPB_SEL_STD;
   input EXE_MEM_WR;
   input MEM_WB_WR;
   output [2:0] MUX_OPA_SEL;
   output [2:0] MUX_OPB_SEL;

   // Internal wires
   wire n25;
   wire n26;
   wire n27;
   wire n28;
   wire n29;
   wire n30;
   wire n31;
   wire n32;
   wire n33;
   wire n34;
   wire n35;
   wire n36;
   wire n37;
   wire n38;
   wire n40;
   wire n41;
   wire n42;
   wire n43;
   wire n44;
   wire n45;
   wire n46;
   wire n47;
   wire n48;
   wire n49;
   wire n50;
   wire n51;
   wire n52;
   wire n53;
   wire n54;
   wire n55;
   wire n56;
   wire n57;
   wire n58;
   wire n4;
   wire n6;
   wire n7;
   wire n9;
   wire n10;
   wire n15;
   wire n16;
   wire n17;
   wire n18;
   wire n19;
   wire n20;

   XOR2_X1 U41 (.A(RD_EX_MEM[2]),
	.B(RS2_ID_EX[2]),
	.Z(n34));
   XOR2_X1 U42 (.A(RD_EX_MEM[0]),
	.B(RS2_ID_EX[0]),
	.Z(n33));
   XOR2_X1 U43 (.A(RD_MEM_WB[2]),
	.B(RS2_ID_EX[2]),
	.Z(n41));
   XOR2_X1 U44 (.A(RD_MEM_WB[0]),
	.B(RS2_ID_EX[0]),
	.Z(n40));
   XOR2_X1 U45 (.A(RD_EX_MEM[2]),
	.B(RS1_ID_EX[2]),
	.Z(n50));
   XOR2_X1 U46 (.A(RD_EX_MEM[0]),
	.B(RS1_ID_EX[0]),
	.Z(n49));
   XOR2_X1 U47 (.A(RD_MEM_WB[2]),
	.B(RS1_ID_EX[2]),
	.Z(n57));
   XOR2_X1 U48 (.A(RD_MEM_WB[0]),
	.B(RS1_ID_EX[0]),
	.Z(n56));
   INV_X1 U3 (.A(n42),
	.ZN(MUX_OPA_SEL[2]));
   NOR4_X1 U5 (.A1(n51),
	.A2(RD_EX_MEM[2]),
	.A3(RD_EX_MEM[3]),
	.A4(RD_EX_MEM[4]),
	.ZN(n32));
   NOR4_X1 U9 (.A1(n58),
	.A2(RD_MEM_WB[4]),
	.A3(RD_MEM_WB[2]),
	.A4(RD_MEM_WB[3]),
	.ZN(n4));
   AND3_X1 U11 (.A1(n47),
	.A2(n46),
	.A3(n45),
	.ZN(n6));
   AND2_X1 U12 (.A1(n30),
	.A2(n29),
	.ZN(n7));
   OAI21_X1 U14 (.A(n44),
	.B1(n43),
	.B2(n16),
	.ZN(MUX_OPA_SEL[0]));
   AND3_X1 U15 (.A1(n55),
	.A2(n53),
	.A3(n9),
	.ZN(n43));
   AND2_X1 U16 (.A1(n54),
	.A2(n52),
	.ZN(n9));
   AND2_X1 U17 (.A1(n38),
	.A2(n10),
	.ZN(n26));
   OAI21_X1 U18 (.A(n27),
	.B1(n26),
	.B2(n17),
	.ZN(MUX_OPB_SEL[1]));
   AND3_X1 U19 (.A1(n35),
	.A2(n37),
	.A3(n36),
	.ZN(n10));
   NAND2_X1 U20 (.A1(n6),
	.A2(n48),
	.ZN(n44));
   OAI21_X1 U21 (.A(n44),
	.B1(n43),
	.B2(n15),
	.ZN(MUX_OPA_SEL[1]));
   NAND3_X1 U22 (.A1(n7),
	.A2(n28),
	.A3(n31),
	.ZN(n27));
   INV_X1 U24 (.A(MUX_OPB_SEL_STD[0]),
	.ZN(n18));
   INV_X1 U25 (.A(MUX_OPB_SEL_STD[1]),
	.ZN(n17));
   INV_X1 U26 (.A(MUX_OPA_SEL_STD[1]),
	.ZN(n15));
   INV_X1 U27 (.A(MUX_OPA_SEL_STD[0]),
	.ZN(n16));
   XNOR2_X1 U28 (.A(RD_MEM_WB[4]),
	.B(RS1_ID_EX[4]),
	.ZN(n53));
   XNOR2_X1 U29 (.A(RD_MEM_WB[3]),
	.B(RS1_ID_EX[3]),
	.ZN(n54));
   OAI21_X1 U30 (.A(n44),
	.B1(n43),
	.B2(MUX_OPA_SEL_STD[2]),
	.ZN(n42));
   XNOR2_X1 U31 (.A(RD_MEM_WB[4]),
	.B(RS2_ID_EX[4]),
	.ZN(n35));
   XNOR2_X1 U32 (.A(RD_MEM_WB[3]),
	.B(RS2_ID_EX[3]),
	.ZN(n37));
   INV_X1 U33 (.A(MEM_WB_WR),
	.ZN(n20));
   INV_X1 U34 (.A(EXE_MEM_WR),
	.ZN(n19));
   OAI21_X1 U35 (.A(n27),
	.B1(n18),
	.B2(n26),
	.ZN(MUX_OPB_SEL[0]));
   NOR4_X1 U36 (.A1(n32),
	.A2(n19),
	.A3(n49),
	.A4(n50),
	.ZN(n48));
   XNOR2_X1 U37 (.A(RD_EX_MEM[3]),
	.B(RS2_ID_EX[3]),
	.ZN(n30));
   XNOR2_X1 U38 (.A(RD_EX_MEM[3]),
	.B(RS1_ID_EX[3]),
	.ZN(n47));
   XNOR2_X1 U39 (.A(RD_EX_MEM[4]),
	.B(RS2_ID_EX[4]),
	.ZN(n28));
   XNOR2_X1 U40 (.A(RD_EX_MEM[4]),
	.B(RS1_ID_EX[4]),
	.ZN(n46));
   OAI21_X1 U49 (.A(n27),
	.B1(n26),
	.B2(MUX_OPB_SEL_STD[2]),
	.ZN(n25));
   XNOR2_X1 U50 (.A(RD_EX_MEM[1]),
	.B(RS2_ID_EX[1]),
	.ZN(n29));
   XNOR2_X1 U51 (.A(RD_EX_MEM[1]),
	.B(RS1_ID_EX[1]),
	.ZN(n45));
   NOR4_X1 U52 (.A1(n32),
	.A2(n33),
	.A3(n34),
	.A4(n19),
	.ZN(n31));
   XNOR2_X1 U53 (.A(RD_MEM_WB[1]),
	.B(RS2_ID_EX[1]),
	.ZN(n36));
   XNOR2_X1 U54 (.A(RD_MEM_WB[1]),
	.B(RS1_ID_EX[1]),
	.ZN(n52));
   OR2_X1 U55 (.A1(RD_EX_MEM[0]),
	.A2(RD_EX_MEM[1]),
	.ZN(n51));
   INV_X1 U56 (.A(n25),
	.ZN(MUX_OPB_SEL[2]));
   NOR4_X1 U57 (.A1(n56),
	.A2(n20),
	.A3(n4),
	.A4(n57),
	.ZN(n55));
   NOR4_X1 U58 (.A1(n40),
	.A2(n4),
	.A3(n41),
	.A4(n20),
	.ZN(n38));
   OR2_X1 U59 (.A1(RD_MEM_WB[1]),
	.A2(RD_MEM_WB[0]),
	.ZN(n58));
endmodule

module FWD_DEC (
	RS1_IF_ID, 
	RS2_IF_ID, 
	IS_COND_JUMP, 
	RD_EX_MEM, 
	RD_MEM_WB, 
	MUX_REGA_SEL, 
	MUX_REGB_SEL);
   input [4:0] RS1_IF_ID;
   input [4:0] RS2_IF_ID;
   input IS_COND_JUMP;
   input [4:0] RD_EX_MEM;
   input [4:0] RD_MEM_WB;
   output [1:0] MUX_REGA_SEL;
   output [1:0] MUX_REGB_SEL;

   // Internal wires
   wire n22;
   wire n23;
   wire n24;
   wire n25;
   wire n26;
   wire n27;
   wire n28;
   wire n29;
   wire n30;
   wire n31;
   wire n32;
   wire n33;
   wire n34;
   wire n35;
   wire n36;
   wire n37;
   wire n38;
   wire n39;
   wire n40;
   wire n41;
   wire n42;
   wire n43;
   wire n44;
   wire n45;
   wire n46;
   wire n47;
   wire n48;
   wire n49;
   wire n50;
   wire n51;
   wire n3;
   wire n4;
   wire n5;

   XOR2_X1 U29 (.A(RS2_IF_ID[1]),
	.B(RD_MEM_WB[1]),
	.Z(n27));
   XOR2_X1 U30 (.A(RS2_IF_ID[4]),
	.B(RD_MEM_WB[4]),
	.Z(n26));
   XOR2_X1 U31 (.A(RS2_IF_ID[3]),
	.B(RD_MEM_WB[3]),
	.Z(n25));
   XOR2_X1 U32 (.A(RS2_IF_ID[2]),
	.B(RD_EX_MEM[2]),
	.Z(n36));
   XOR2_X1 U33 (.A(RS2_IF_ID[0]),
	.B(RD_EX_MEM[0]),
	.Z(n35));
   XOR2_X1 U34 (.A(RS1_IF_ID[1]),
	.B(RD_MEM_WB[1]),
	.Z(n41));
   XOR2_X1 U35 (.A(RS1_IF_ID[4]),
	.B(RD_MEM_WB[4]),
	.Z(n40));
   XOR2_X1 U36 (.A(RS1_IF_ID[3]),
	.B(RD_MEM_WB[3]),
	.Z(n39));
   XOR2_X1 U37 (.A(RS1_IF_ID[2]),
	.B(RD_EX_MEM[2]),
	.Z(n50));
   XOR2_X1 U38 (.A(RS1_IF_ID[0]),
	.B(RD_EX_MEM[0]),
	.Z(n49));
   INV_X1 U2 (.A(IS_COND_JUMP),
	.ZN(n5));
   INV_X1 U3 (.A(n23),
	.ZN(MUX_REGA_SEL[0]));
   INV_X1 U4 (.A(n22),
	.ZN(MUX_REGB_SEL[0]));
   NOR4_X1 U5 (.A1(RS1_IF_ID[3]),
	.A2(RS1_IF_ID[4]),
	.A3(RS1_IF_ID[2]),
	.A4(n51),
	.ZN(n48));
   OR2_X1 U6 (.A1(RS1_IF_ID[1]),
	.A2(RS1_IF_ID[0]),
	.ZN(n51));
   NOR4_X1 U7 (.A1(n38),
	.A2(n39),
	.A3(n40),
	.A4(n41),
	.ZN(MUX_REGA_SEL[1]));
   NOR4_X1 U8 (.A1(n24),
	.A2(n25),
	.A3(n26),
	.A4(n27),
	.ZN(MUX_REGB_SEL[1]));
   NOR4_X1 U9 (.A1(n48),
	.A2(n5),
	.A3(n49),
	.A4(n50),
	.ZN(n47));
   NOR4_X1 U10 (.A1(n34),
	.A2(n5),
	.A3(n35),
	.A4(n36),
	.ZN(n33));
   NAND4_X1 U11 (.A1(n44),
	.A2(n45),
	.A3(n46),
	.A4(n47),
	.ZN(n23));
   NAND4_X1 U12 (.A1(n30),
	.A2(n31),
	.A3(n32),
	.A4(n33),
	.ZN(n22));
   NAND4_X1 U13 (.A1(n42),
	.A2(n43),
	.A3(n4),
	.A4(n23),
	.ZN(n38));
   XNOR2_X1 U14 (.A(RD_MEM_WB[2]),
	.B(RS1_IF_ID[2]),
	.ZN(n42));
   INV_X1 U15 (.A(n48),
	.ZN(n4));
   NAND4_X1 U16 (.A1(n28),
	.A2(n29),
	.A3(n3),
	.A4(n22),
	.ZN(n24));
   XNOR2_X1 U17 (.A(RD_MEM_WB[2]),
	.B(RS2_IF_ID[2]),
	.ZN(n28));
   INV_X1 U18 (.A(n34),
	.ZN(n3));
   NOR4_X1 U19 (.A1(RS2_IF_ID[3]),
	.A2(RS2_IF_ID[4]),
	.A3(RS2_IF_ID[2]),
	.A4(n37),
	.ZN(n34));
   OR2_X1 U20 (.A1(RS2_IF_ID[1]),
	.A2(RS2_IF_ID[0]),
	.ZN(n37));
   XNOR2_X1 U21 (.A(RD_EX_MEM[3]),
	.B(RS1_IF_ID[3]),
	.ZN(n46));
   XNOR2_X1 U22 (.A(RD_EX_MEM[3]),
	.B(RS2_IF_ID[3]),
	.ZN(n32));
   XNOR2_X1 U23 (.A(RD_EX_MEM[4]),
	.B(RS1_IF_ID[4]),
	.ZN(n45));
   XNOR2_X1 U24 (.A(RD_EX_MEM[4]),
	.B(RS2_IF_ID[4]),
	.ZN(n30));
   XNOR2_X1 U25 (.A(RD_EX_MEM[1]),
	.B(RS1_IF_ID[1]),
	.ZN(n44));
   XNOR2_X1 U26 (.A(RD_EX_MEM[1]),
	.B(RS2_IF_ID[1]),
	.ZN(n31));
   XNOR2_X1 U27 (.A(RD_MEM_WB[0]),
	.B(RS2_IF_ID[0]),
	.ZN(n29));
   XNOR2_X1 U28 (.A(RD_MEM_WB[0]),
	.B(RS1_IF_ID[0]),
	.ZN(n43));
endmodule

module HDU (
	RS1_IF_ID, 
	RS2_IF_ID, 
	RD_ID_EXE, 
	RD_EXE_MEM, 
	MEM_LD_EXE, 
	MEM_LD_MEM, 
	IS_COND_JUMP, 
	STALL);
   input [4:0] RS1_IF_ID;
   input [4:0] RS2_IF_ID;
   input [4:0] RD_ID_EXE;
   input [4:0] RD_EXE_MEM;
   input MEM_LD_EXE;
   input MEM_LD_MEM;
   input IS_COND_JUMP;
   output STALL;

   // Internal wires
   wire n18;
   wire n19;
   wire n20;
   wire n21;
   wire n22;
   wire n23;
   wire n24;
   wire n25;
   wire n26;
   wire n27;
   wire n28;
   wire n29;
   wire n30;
   wire n31;
   wire n32;
   wire n33;
   wire n34;
   wire n35;
   wire n36;
   wire n37;
   wire n38;
   wire n39;
   wire n40;
   wire n41;
   wire n42;
   wire n43;
   wire n44;
   wire n45;
   wire n1;

   OAI33_X1 U18 (.A1(n22),
	.A2(n23),
	.A3(n24),
	.B1(n25),
	.B2(n26),
	.B3(n27),
	.ZN(n20));
   XOR2_X1 U19 (.A(RS2_IF_ID[4]),
	.B(RD_ID_EXE[4]),
	.Z(n27));
   XOR2_X1 U20 (.A(RS2_IF_ID[3]),
	.B(RD_ID_EXE[3]),
	.Z(n26));
   NAND3_X1 U21 (.A1(n28),
	.A2(n29),
	.A3(n30),
	.ZN(n25));
   XOR2_X1 U22 (.A(RS1_IF_ID[4]),
	.B(RD_ID_EXE[4]),
	.Z(n24));
   XOR2_X1 U23 (.A(RS1_IF_ID[3]),
	.B(RD_ID_EXE[3]),
	.Z(n23));
   NAND3_X1 U24 (.A1(n31),
	.A2(n32),
	.A3(n33),
	.ZN(n22));
   OAI33_X1 U25 (.A1(n34),
	.A2(n35),
	.A3(n36),
	.B1(n37),
	.B2(n38),
	.B3(n39),
	.ZN(n21));
   XOR2_X1 U26 (.A(RS2_IF_ID[4]),
	.B(RD_EXE_MEM[4]),
	.Z(n39));
   XOR2_X1 U27 (.A(RS2_IF_ID[3]),
	.B(RD_EXE_MEM[3]),
	.Z(n38));
   NAND3_X1 U28 (.A1(n40),
	.A2(n41),
	.A3(n42),
	.ZN(n37));
   XOR2_X1 U29 (.A(RS1_IF_ID[4]),
	.B(RD_EXE_MEM[4]),
	.Z(n36));
   XOR2_X1 U30 (.A(RS1_IF_ID[3]),
	.B(RD_EXE_MEM[3]),
	.Z(n35));
   NAND3_X1 U31 (.A1(n43),
	.A2(n44),
	.A3(n45),
	.ZN(n34));
   OAI21_X1 U2 (.A(n19),
	.B1(n18),
	.B2(n1),
	.ZN(STALL));
   INV_X1 U3 (.A(IS_COND_JUMP),
	.ZN(n1));
   NAND2_X1 U4 (.A1(MEM_LD_EXE),
	.A2(n20),
	.ZN(n19));
   AOI21_X1 U5 (.A(n20),
	.B1(MEM_LD_MEM),
	.B2(n21),
	.ZN(n18));
   XNOR2_X1 U6 (.A(RD_ID_EXE[1]),
	.B(RS2_IF_ID[1]),
	.ZN(n29));
   XNOR2_X1 U7 (.A(RD_ID_EXE[0]),
	.B(RS2_IF_ID[0]),
	.ZN(n28));
   XNOR2_X1 U8 (.A(RD_ID_EXE[2]),
	.B(RS2_IF_ID[2]),
	.ZN(n30));
   XNOR2_X1 U9 (.A(RD_ID_EXE[1]),
	.B(RS1_IF_ID[1]),
	.ZN(n32));
   XNOR2_X1 U10 (.A(RD_ID_EXE[0]),
	.B(RS1_IF_ID[0]),
	.ZN(n31));
   XNOR2_X1 U11 (.A(RD_ID_EXE[2]),
	.B(RS1_IF_ID[2]),
	.ZN(n33));
   XNOR2_X1 U12 (.A(RD_EXE_MEM[0]),
	.B(RS2_IF_ID[0]),
	.ZN(n40));
   XNOR2_X1 U13 (.A(RD_EXE_MEM[0]),
	.B(RS1_IF_ID[0]),
	.ZN(n43));
   XNOR2_X1 U14 (.A(RD_EXE_MEM[2]),
	.B(RS1_IF_ID[2]),
	.ZN(n45));
   XNOR2_X1 U15 (.A(RD_EXE_MEM[2]),
	.B(RS2_IF_ID[2]),
	.ZN(n42));
   XNOR2_X1 U16 (.A(RD_EXE_MEM[1]),
	.B(RS2_IF_ID[1]),
	.ZN(n41));
   XNOR2_X1 U17 (.A(RD_EXE_MEM[1]),
	.B(RS1_IF_ID[1]),
	.ZN(n44));
endmodule

module CU (
	clk, 
	rst, 
	OPCODE, 
	FUNC3, 
	EQU, 
	RS1_IF_ID, 
	RS2_IF_ID, 
	RS1_ID_EXE, 
	RS2_ID_EXE, 
	RD_ID_EXE, 
	RD_EXE_MEM, 
	RD_MEM_WB, 
	DRAM_WR_IN, 
	DRAM_RD_IN, 
	DRAM_EN, 
	RF_RD1, 
	RF_RD2, 
	RF_WR, 
	JUMP, 
	MUX_SEL_WB, 
	FETCH_EN, 
	DECODE_EN, 
	EXE_EN, 
	MEM_EN, 
	WB_EN, 
	RF_OUT1_SEL, 
	RF_OUT2_SEL, 
	ALU_OPA_SEL, 
	ALU_OPB_SEL, 
	MUX_SEL_IMM, 
	ALU_OP);
   input clk;
   input rst;
   input [6:0] OPCODE;
   input [2:0] FUNC3;
   input EQU;
   input [4:0] RS1_IF_ID;
   input [4:0] RS2_IF_ID;
   input [4:0] RS1_ID_EXE;
   input [4:0] RS2_ID_EXE;
   input [4:0] RD_ID_EXE;
   input [4:0] RD_EXE_MEM;
   input [4:0] RD_MEM_WB;
   output DRAM_WR_IN;
   output DRAM_RD_IN;
   output DRAM_EN;
   output RF_RD1;
   output RF_RD2;
   output RF_WR;
   output JUMP;
   output MUX_SEL_WB;
   output FETCH_EN;
   output DECODE_EN;
   output EXE_EN;
   output MEM_EN;
   output WB_EN;
   output [1:0] RF_OUT1_SEL;
   output [1:0] RF_OUT2_SEL;
   output [2:0] ALU_OPA_SEL;
   output [2:0] ALU_OPB_SEL;
   output [2:0] MUX_SEL_IMM;
   output [2:0] ALU_OP;

   // Internal wires
   wire FE_PHN139_n13;
   wire FE_PHN138_n8;
   wire FE_PHN137_n16;
   wire IS_COND_JUMP;
   wire ctrl_word_E_3_;
   wire ctrl_word_M_0_;
   wire STALL;
   wire N98;
   wire N99;
   wire N102;
   wire N104;
   wire N105;
   wire N106;
   wire N107;
   wire N108;
   wire N112;
   wire N117;
   wire N118;
   wire N119;
   wire n4;
   wire n6;
   wire n8;
   wire n13;
   wire n14;
   wire n16;
   wire n17;
   wire n36;
   wire n37;
   wire n38;
   wire n39;
   wire n40;
   wire n41;
   wire n42;
   wire n43;
   wire n44;
   wire n45;
   wire n46;
   wire n47;
   wire n48;
   wire n49;
   wire n50;
   wire n51;
   wire n52;
   wire n53;
   wire n54;
   wire n55;
   wire n56;
   wire n57;
   wire n5;
   wire n7;
   wire n9;
   wire n11;
   wire n15;
   wire n18;
   wire n19;
   wire n20;
   wire n21;
   wire n22;
   wire n23;
   wire n26;
   wire n28;
   wire n29;
   wire n34;
   wire n58;
   wire n59;
   wire n60;
   wire n61;
   wire n62;
   wire n64;
   wire n65;
   wire n66;
   wire n67;
   wire n68;
   wire n69;
   wire n70;
   wire [2:0] MUX_OPA_SEL_STD;
   wire [2:0] MUX_OPB_SEL_STD;

   assign DECODE_EN = FETCH_EN ;

   BUF_X1 FE_PHC139_n13 (.A(n13),
	.Z(FE_PHN139_n13));
   BUF_X1 FE_PHC138_n8 (.A(n8),
	.Z(FE_PHN138_n8));
   BUF_X1 FE_PHC137_n16 (.A(n16),
	.Z(FE_PHN137_n16));
   DFF_X1 alu_ctrl1_reg_2_ (.D(N119),
	.CK(clk),
	.Q(ALU_OP[2]));
   DFF_X1 alu_ctrl1_reg_1_ (.D(N118),
	.CK(clk),
	.Q(ALU_OP[1]));
   DFF_X1 alu_ctrl1_reg_0_ (.D(N117),
	.CK(clk),
	.Q(ALU_OP[0]));
   DFF_X1 ctrl_word_M_reg_3_ (.D(N112),
	.CK(clk),
	.Q(DRAM_RD_IN));
   DFF_X1 ctrl_word_E_reg_0_ (.D(N98),
	.CK(clk),
	.QN(n17));
   DFF_X1 ctrl_word_E_reg_11_ (.D(N108),
	.CK(clk),
	.Q(MUX_OPA_SEL_STD[1]));
   DFF_X1 ctrl_word_E_reg_10_ (.D(N107),
	.CK(clk),
	.Q(MUX_OPA_SEL_STD[0]));
   DFF_X1 ctrl_word_E_reg_8_ (.D(N106),
	.CK(clk),
	.Q(MUX_OPB_SEL_STD[1]));
   DFF_X1 ctrl_word_E_reg_4_ (.D(N102),
	.CK(clk),
	.QN(n16));
   DFF_X1 ctrl_word_E_reg_7_ (.D(N105),
	.CK(clk),
	.Q(MUX_OPB_SEL_STD[0]));
   DFF_X1 ctrl_word_E_reg_1_ (.D(N99),
	.CK(clk),
	.QN(n14));
   DFF_X1 ctrl_word_E_reg_3_ (.D(N99),
	.CK(clk),
	.Q(ctrl_word_E_3_));
   DFF_X1 ctrl_word_E_reg_6_ (.D(N104),
	.CK(clk),
	.Q(MEM_EN));
   DFF_X1 ctrl_word_E_reg_2_ (.D(N104),
	.CK(clk),
	.QN(n8));
   NAND3_X1 U72 (.A1(IS_COND_JUMP),
	.A2(FETCH_EN),
	.A3(EQU),
	.ZN(n52));
   FWD_EXE forward_unit_exe (.RS1_ID_EX(RS1_ID_EXE),
	.RS2_ID_EX(RS2_ID_EXE),
	.RD_EX_MEM(RD_EXE_MEM),
	.RD_MEM_WB(RD_MEM_WB),
	.MUX_OPA_SEL_STD({ 1'b0,
		MUX_OPA_SEL_STD[1],
		MUX_OPA_SEL_STD[0] }),
	.MUX_OPB_SEL_STD({ 1'b0,
		MUX_OPB_SEL_STD[1],
		MUX_OPB_SEL_STD[0] }),
	.EXE_MEM_WR(ctrl_word_M_0_),
	.MEM_WB_WR(RF_WR),
	.MUX_OPA_SEL(ALU_OPA_SEL),
	.MUX_OPB_SEL(ALU_OPB_SEL));
   FWD_DEC forward_unit_dec (.RS1_IF_ID(RS1_IF_ID),
	.RS2_IF_ID(RS2_IF_ID),
	.IS_COND_JUMP(IS_COND_JUMP),
	.RD_EX_MEM(RD_EXE_MEM),
	.RD_MEM_WB(RD_MEM_WB),
	.MUX_REGA_SEL(RF_OUT1_SEL),
	.MUX_REGB_SEL(RF_OUT2_SEL));
   HDU hazard_unit (.RS1_IF_ID(RS1_IF_ID),
	.RS2_IF_ID(RS2_IF_ID),
	.RD_ID_EXE(RD_ID_EXE),
	.RD_EXE_MEM(RD_EXE_MEM),
	.MEM_LD_EXE(ctrl_word_E_3_),
	.MEM_LD_MEM(DRAM_RD_IN),
	.IS_COND_JUMP(IS_COND_JUMP),
	.STALL(STALL));
   DFF_X1 ctrl_word_W_reg_1_ (.D(n22),
	.CK(clk),
	.Q(MUX_SEL_WB));
   DFF_X1 ctrl_word_W_reg_0_ (.D(n21),
	.CK(clk),
	.Q(RF_WR));
   DFF_X1 ctrl_word_M_reg_5_ (.D(n20),
	.CK(clk),
	.Q(DRAM_EN));
   DFF_X1 ctrl_word_M_reg_4_ (.D(n19),
	.CK(clk),
	.Q(DRAM_WR_IN));
   DFF_X1 ctrl_word_M_reg_2_ (.D(n18),
	.CK(clk),
	.Q(WB_EN));
   DFF_X1 ctrl_word_M_reg_0_ (.D(n15),
	.CK(clk),
	.Q(ctrl_word_M_0_),
	.QN(n4));
   DFF_X1 ctrl_word_M_reg_1_ (.D(n11),
	.CK(clk),
	.QN(n6));
   DFF_X1 ctrl_word_E_reg_5_ (.D(n9),
	.CK(clk),
	.QN(n13));
   OR2_X1 U5 (.A1(n47),
	.A2(n7),
	.ZN(n26));
   AND2_X1 U7 (.A1(OPCODE[1]),
	.A2(OPCODE[6]),
	.ZN(n5));
   OR2_X1 U8 (.A1(n66),
	.A2(OPCODE[2]),
	.ZN(n7));
   NOR2_X1 U9 (.A1(n60),
	.A2(n41),
	.ZN(n9));
   NOR2_X1 U10 (.A1(n14),
	.A2(rst),
	.ZN(n11));
   NOR2_X1 U12 (.A1(n17),
	.A2(rst),
	.ZN(n15));
   NOR2_X1 U16 (.A1(FE_PHN138_n8),
	.A2(rst),
	.ZN(n18));
   NOR2_X1 U17 (.A1(FE_PHN137_n16),
	.A2(rst),
	.ZN(n19));
   NOR2_X1 U18 (.A1(FE_PHN139_n13),
	.A2(rst),
	.ZN(n20));
   NOR2_X1 U19 (.A1(n4),
	.A2(rst),
	.ZN(n21));
   NOR2_X1 U20 (.A1(n6),
	.A2(rst),
	.ZN(n22));
   INV_X1 U21 (.A(n26),
	.ZN(n42));
   AND3_X1 U22 (.A1(n55),
	.A2(OPCODE[5]),
	.A3(n5),
	.ZN(n23));
   AND2_X1 U23 (.A1(n57),
	.A2(n28),
	.ZN(n56));
   NAND3_X1 U26 (.A1(n55),
	.A2(OPCODE[5]),
	.A3(n5),
	.ZN(n54));
   NOR3_X1 U28 (.A1(OPCODE[2]),
	.A2(OPCODE[3]),
	.A3(n54),
	.ZN(IS_COND_JUMP));
   INV_X1 U29 (.A(n29),
	.ZN(n48));
   NOR2_X1 U30 (.A1(OPCODE[2]),
	.A2(OPCODE[4]),
	.ZN(n28));
   AND3_X1 U31 (.A1(OPCODE[2]),
	.A2(n23),
	.A3(OPCODE[3]),
	.ZN(n29));
   AND2_X1 U32 (.A1(n37),
	.A2(n64),
	.ZN(n40));
   NAND2_X1 U33 (.A1(n51),
	.A2(n26),
	.ZN(MUX_SEL_IMM[1]));
   AND2_X1 U34 (.A1(n49),
	.A2(n65),
	.ZN(n37));
   INV_X1 U35 (.A(n38),
	.ZN(n62));
   NAND4_X1 U36 (.A1(n49),
	.A2(n64),
	.A3(n65),
	.A4(n53),
	.ZN(EXE_EN));
   AND2_X1 U37 (.A1(n62),
	.A2(n51),
	.ZN(n53));
   AOI21_X1 U38 (.A(n41),
	.B1(n37),
	.B2(n62),
	.ZN(N107));
   NOR2_X1 U39 (.A1(n41),
	.A2(n61),
	.ZN(N104));
   INV_X1 U40 (.A(EXE_EN),
	.ZN(n61));
   NOR2_X1 U41 (.A1(n41),
	.A2(n49),
	.ZN(N99));
   INV_X1 U42 (.A(MUX_SEL_IMM[2]),
	.ZN(n64));
   OAI21_X1 U43 (.A(n34),
	.B1(n40),
	.B2(n41),
	.ZN(N105));
   INV_X1 U44 (.A(N102),
	.ZN(n34));
   NOR2_X1 U45 (.A1(n67),
	.A2(n47),
	.ZN(MUX_SEL_IMM[2]));
   NAND2_X1 U46 (.A1(n50),
	.A2(n48),
	.ZN(MUX_SEL_IMM[0]));
   NOR2_X1 U47 (.A1(IS_COND_JUMP),
	.A2(n29),
	.ZN(n51));
   NAND2_X1 U48 (.A1(n52),
	.A2(n48),
	.ZN(JUMP));
   NOR2_X1 U49 (.A1(n38),
	.A2(IS_COND_JUMP),
	.ZN(n36));
   NAND2_X1 U50 (.A1(n56),
	.A2(n66),
	.ZN(n49));
   NAND2_X1 U51 (.A1(n26),
	.A2(n50),
	.ZN(n38));
   INV_X1 U52 (.A(n46),
	.ZN(n65));
   NAND2_X1 U53 (.A1(n37),
	.A2(n36),
	.ZN(RF_RD1));
   INV_X1 U54 (.A(n36),
	.ZN(RF_RD2));
   NAND2_X1 U55 (.A1(FETCH_EN),
	.A2(n70),
	.ZN(n41));
   NOR4_X1 U56 (.A1(n66),
	.A2(n47),
	.A3(n41),
	.A4(n67),
	.ZN(N108));
   NOR2_X1 U57 (.A1(n50),
	.A2(n41),
	.ZN(N102));
   AOI21_X1 U58 (.A(n41),
	.B1(n39),
	.B2(n40),
	.ZN(N98));
   NOR2_X1 U59 (.A1(n29),
	.A2(n42),
	.ZN(n39));
   NAND2_X1 U60 (.A1(n42),
	.A2(n59),
	.ZN(n43));
   NOR2_X1 U61 (.A1(n41),
	.A2(n48),
	.ZN(N106));
   INV_X1 U62 (.A(n56),
	.ZN(n60));
   NOR4_X1 U63 (.A1(n68),
	.A2(n69),
	.A3(OPCODE[3]),
	.A4(OPCODE[6]),
	.ZN(n57));
   INV_X1 U64 (.A(OPCODE[1]),
	.ZN(n68));
   NOR2_X1 U65 (.A1(OPCODE[4]),
	.A2(n69),
	.ZN(n55));
   NAND2_X1 U66 (.A1(OPCODE[4]),
	.A2(n57),
	.ZN(n47));
   NAND2_X1 U67 (.A1(n56),
	.A2(OPCODE[5]),
	.ZN(n50));
   INV_X1 U68 (.A(OPCODE[5]),
	.ZN(n66));
   INV_X1 U69 (.A(OPCODE[2]),
	.ZN(n67));
   NOR3_X1 U70 (.A1(OPCODE[2]),
	.A2(OPCODE[5]),
	.A3(n47),
	.ZN(n46));
   INV_X1 U71 (.A(STALL),
	.ZN(FETCH_EN));
   OAI21_X1 U73 (.A(n70),
	.B1(FUNC3[2]),
	.B2(FUNC3[1]),
	.ZN(n44));
   NOR4_X1 U74 (.A1(n44),
	.A2(n65),
	.A3(n59),
	.A4(n58),
	.ZN(N117));
   INV_X1 U75 (.A(FUNC3[2]),
	.ZN(n58));
   AOI211_X1 U76 (.A(n44),
	.B(FUNC3[1]),
	.C1(n43),
	.C2(n45),
	.ZN(N118));
   NAND2_X1 U77 (.A1(FUNC3[0]),
	.A2(n46),
	.ZN(n45));
   INV_X1 U78 (.A(rst),
	.ZN(n70));
   NOR3_X1 U79 (.A1(n43),
	.A2(FUNC3[2]),
	.A3(n44),
	.ZN(N119));
   INV_X1 U80 (.A(FUNC3[0]),
	.ZN(n59));
   AND2_X1 U81 (.A1(ctrl_word_E_3_),
	.A2(n70),
	.ZN(N112));
   INV_X1 U82 (.A(OPCODE[0]),
	.ZN(n69));
endmodule

module RISCV (
	clk, 
	rst, 
	en, 
	IRAM_OUT, 
	DRAM_OUT, 
	IRAM_ADDR, 
	DRAM_EN, 
	DRAM_IN, 
	DRAM_ADDR, 
	DRAM_WR, 
	DRAM_RD);
   input clk;
   input rst;
   input en;
   input [31:0] IRAM_OUT;
   input [31:0] DRAM_OUT;
   output [31:0] IRAM_ADDR;
   output DRAM_EN;
   output [31:0] DRAM_IN;
   output [31:0] DRAM_ADDR;
   output DRAM_WR;
   output DRAM_RD;

   // Internal wires
   wire FETCH_EN_c;
   wire DECODE_EN_c;
   wire EXE_EN_c;
   wire MEM_EN_c;
   wire WB_EN_c;
   wire DRAM_WR_IN_c;
   wire DRAM_RD_IN_c;
   wire RF_RD1_c;
   wire RF_RD2_c;
   wire RF_WR_c;
   wire JUMP_c;
   wire MUX_SEL_WB_c;
   wire EQU_s;
   wire [1:0] RF_OUT1_SEL;
   wire [1:0] RF_OUT2_SEL;
   wire [2:0] ALU_OPA_SEL_c;
   wire [2:0] ALU_OPB_SEL_c;
   wire [2:0] MUX_SEL_IMM_c;
   wire [2:0] ALU_OP_c;
   wire [6:0] OPCODE_s;
   wire [2:0] FUNC3_s;
   wire [4:0] RS1_IF_ID;
   wire [4:0] RS2_IF_ID;
   wire [4:0] RS1_ID_EXE;
   wire [4:0] RS2_ID_EXE;
   wire [4:0] RD_EXE_MEM;
   wire [4:0] RD_MEM_WB;
   wire [4:0] RD_ID_EXE;

   DP DP_u (.clk(clk),
	.rst(rst),
	.FETCH_EN(FETCH_EN_c),
	.DECODE_EN(DECODE_EN_c),
	.EXE_EN(EXE_EN_c),
	.MEM_EN(MEM_EN_c),
	.WB_EN(WB_EN_c),
	.IRAM_OUT(IRAM_OUT),
	.DRAM_OUT(DRAM_OUT),
	.DRAM_WR_IN(DRAM_WR_IN_c),
	.DRAM_RD_IN(DRAM_RD_IN_c),
	.RF_RD1(RF_RD1_c),
	.RF_RD2(RF_RD2_c),
	.RF_WR(RF_WR_c),
	.JUMP(JUMP_c),
	.MUX_SEL_WB(MUX_SEL_WB_c),
	.RF_OUT1_SEL(RF_OUT1_SEL),
	.RF_OUT2_SEL(RF_OUT2_SEL),
	.ALU_OPA_SEL(ALU_OPA_SEL_c),
	.ALU_OPB_SEL(ALU_OPB_SEL_c),
	.MUX_SEL_IMM(MUX_SEL_IMM_c),
	.ALU_OP(ALU_OP_c),
	.IRAM_ADDR(IRAM_ADDR),
	.DRAM_IN(DRAM_IN),
	.DRAM_ADDR(DRAM_ADDR),
	.DRAM_WR(DRAM_WR),
	.DRAM_RD(DRAM_RD),
	.OPCODE(OPCODE_s),
	.FUNC3(FUNC3_s),
	.EQU(EQU_s),
	.RS1_IF_ID(RS1_IF_ID),
	.RS2_IF_ID(RS2_IF_ID),
	.RS1_ID_EXE(RS1_ID_EXE),
	.RS2_ID_EXE(RS2_ID_EXE),
	.RD_EXE_MEM(RD_EXE_MEM),
	.RD_MEM_WB(RD_MEM_WB),
	.RD_ID_EXE(RD_ID_EXE));
   CU CU_u (.clk(clk),
	.rst(rst),
	.OPCODE(OPCODE_s),
	.FUNC3(FUNC3_s),
	.EQU(EQU_s),
	.RS1_IF_ID(RS1_IF_ID),
	.RS2_IF_ID(RS2_IF_ID),
	.RS1_ID_EXE(RS1_ID_EXE),
	.RS2_ID_EXE(RS2_ID_EXE),
	.RD_ID_EXE(RD_ID_EXE),
	.RD_EXE_MEM(RD_EXE_MEM),
	.RD_MEM_WB(RD_MEM_WB),
	.DRAM_WR_IN(DRAM_WR_IN_c),
	.DRAM_RD_IN(DRAM_RD_IN_c),
	.DRAM_EN(DRAM_EN),
	.RF_RD1(RF_RD1_c),
	.RF_RD2(RF_RD2_c),
	.RF_WR(RF_WR_c),
	.JUMP(JUMP_c),
	.MUX_SEL_WB(MUX_SEL_WB_c),
	.FETCH_EN(FETCH_EN_c),
	.DECODE_EN(DECODE_EN_c),
	.EXE_EN(EXE_EN_c),
	.MEM_EN(MEM_EN_c),
	.WB_EN(WB_EN_c),
	.RF_OUT1_SEL(RF_OUT1_SEL),
	.RF_OUT2_SEL(RF_OUT2_SEL),
	.ALU_OPA_SEL(ALU_OPA_SEL_c),
	.ALU_OPB_SEL(ALU_OPB_SEL_c),
	.MUX_SEL_IMM(MUX_SEL_IMM_c),
	.ALU_OP(ALU_OP_c));
endmodule

